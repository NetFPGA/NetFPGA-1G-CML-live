XlxV64EB    159f     840"b��ҁXc�D�x�۽A$l�e}I��Y���E��_(����N��H�9�7l���+�J9���-:|ǙJTݭR��bP�/9sS�$���^A�v �Y���+�b�<;�ͮ��=3�� ߇��N��Q$n}�E�B4#g�\A4���oW��L��՜��_�Qۜy_\^�� S��W��LOʽTzdgb����E����I-�[�[F#Jv���3lc��c�y͎�T�x�r!�lw�ʦf�'/�F8��R��R#�sb���2��`T��N���qg��)��_l��wd^M��u����ad>�+����\B*��[�wW��[���T2�tӍDk>�ݏ�1�Y�����B����/C�~! A���Q�}�bҕ���XKꞃ<�S��X�̎��g�rK��P����6j�+�q�<\I}K�F�	�����͎���!$]i�\��i:j(��n�On����јo[�
��w�#Y )Qw.\�9�]aGA=f8���T6��H7x^�O?	�����Ьɇ젻O��-o���ytt�����b��'�~��IVQC�F�����A��ז�q?Xx	vb�y�����dc�6;��h��
���jĉ+~�S����J����
�#��㶔;˃�-�~
fa�F�܂���S0�?��)���M���VɡCP��K��e�s�C�,V
K�G�=��i���=����+05DM���cJ¸��O����Σ�h�!�����68.�҆�@6ӥB�1W|m<1�����S���J�
G�����*�[����� �ZH�z�<���
���h+-�Q?�mo����u63��\v�`L����F���Y#YMR|�b��8bA5cb5�e�N}ן[@�`��G�I�pt�z?._����ۜ������dt��I۾>X`���*�x�c�\$���5���1�_n(��Is��m%���{���E"P����\aG �Ÿ��9U���Q1+�C@E]*=�v�8 �]��^�2F*��'���JAB>(�y��j�U�ѴV|��=�l�g-�X�הh�1*����&�'d�~a+�� �A��@/���72�E��G;gKڒ��2�e�V�� �	J2] ���9��@\N��G�n�6u����?!�_G��Gw��򙟰E+�j��м3��8p�?ʉ��픗�w�S��3���w�"3@#D@$sx=�'\"�6�M߂w_~�N���P���`�����Y��#7!��[�L[a�7��8���L)?j��7��P��0ȼA_Hl�Z|OkA�z
�-��9cXܫ���;�j�X���&�d���+ۻ,�k��ӎ��zhZ�=NT��)�=V�h�n��A6�f��Oz���Μ����Z�5����݂�Zr(�}����Gtd�%����c�1{�g}\ň�	���m�|���т���:�7Z6���=��p�Ƅ&�h%�y0�l����O00�V����j�M��sa�!r�<#E��
�_���X�\�z�&�ݤ>Q����:l#QsJ���
e9��m��5��G��9��Tq�YZ�$���@J��c����9���U���9=���ѓXTo�4
h�����c9��iŝb�Z&��ǀ����5�*Zf�_zj�����ĕɺ��N�f�:jt+uDu9�EI	,����f�	���~r��g"?�$T��̬(:����o9��%L��F�T�p���+,/
��-~3l$o�����z7l��T`"�NʆF��/i�/����~&��2>{���GZ2��R�0�����*���F��q�|: �v��S��L`9�#�ٺ>�p7����;��C]��p�8[Za���M_FP����mx\J�r�}-�~�4�s(��ݑ4�Nͫ	-X�P����t��ͫ�5%��	��ƣ@Xqӯ��RX��V�j9�4��ǝ�l뱦�*4\�y�7�,�c�����E*	"!N~3bQCP0G���x�$O�@�7j�.��Uu�9H���l~�e������K���@M��WwrzD��au�\��HG� �|��Ժ�"/����