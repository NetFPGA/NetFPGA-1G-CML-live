XlxV64EB    5d01    10d0�Z5Lo�X�]�dZY�A�TLCr�j1�<�u�rI:��p����9R��c��Ѐ�5$�L-%��&˔¬X��YM�	��f�NY���#*/��]�U+j]�GJ�^.6�]3��ZNߵ��&�ٸ���H�}��<�S�nh�No��R��Y=�;pl!��r{����K�.	k� N`x���9�[���ԓCسu%��R���߈&��1��!��؝q4�?���/㪼F}��+�K�5�?��Z5H�6Mm�������Q�ix�l\���I)����T���̿Fcϧ�� #���ɸ�8�Eʰ�|��!���Xw����_o�?�B��J��S���y���P��)-DS�=f��&�ui{��vk�SP�1_h�
j2�VZ�/{X�be9�k3)Y�A�H=({0hތ���C�g�ڦu���PN����������I�x�%Cn����4��=]��:���LT.�%:?���l4>�
�x�U²�*	�!�3�j����J �'$���+5=�s!���/F�9�oY >�18�?��َ�@�S�#�4�q���QM]Ҽ�?°[�J;�\�+ǎ�~;µ���ln��HZ*U;�1�J~-���Cj��E��&nJ޾�ߨѧ�������Pv�|���Q�[�ܦ��d�)D^�H� 5o���J5�/q@T2ZQ�nН��R��Z��(���vb�|�l7�F�[T<�, 
A�-
(�-������0��0��
ޛ~��"E����P]�ϓ�����8IC�y��J���0�h����P)i��ʍ,�"��/ɉ�%�N����LT��n�Od�&���0��j�Ep	0"���m�ݻ�ԗ�Ϊ2�>2����c�W�f���IXq�]�q_?�-RIJRh��4 ���g]:�Ffg6��5��"-�K�"DZ�ڵ^��������BMns�C�R�0��_A�g�"!�`P���ɯc(�����i.����y���w~֯��o��v�S��UՄ�9i0v�ވ3ɹLD�|}����,���*��=�e���`��nH��yG�Y��K�s�Z9�׮ڥ3�5�ּ�G#���!���0k�19��J�8)b��'���p?�|V??.��!�Uʛ��Ա��7���k��k>p;�юJhU[D���� i�H���
��B	P��0�����y�@Z��Mk\�,8De�Ss��A�C��Zc��D�A^��\�q.[̰�
W��T�0�/��.(��_�\��;�A�j�8�*ਦ���ujS���9�;l5��jq$�6ּ�p����N�^�0�{�L0���e�Ll�s��n���1v�*�@��9�nx+GW�,d��	&��U(��䂛t	�.���1�`��$�c�/F~Y
�Hy_����Q�]
n�xU{�t�+�g>/ٺ��܇����Ŀ~�s�5�Q��Т}�g����tq^}�W������"���iK��,مS�!�In`ʾ��������zP�/rL@��*\t�O���#�SW��6�@Mh�E����c�<H9\������P{�^������^p+OΦ�k���^�ZԤ��(t�J�֜�1y,!\c��#Ӎ��6z�O�W�Є�J\�����/[&�M0:-�UXڶhw�Ra�H�GrL/ݽ�� ��]_�K���4{����ϳf�Y!8��J���X����{�P��Kx�-Ӹ��|qh� @�
#ȉ������>`-��L�N"�[�z�Z�Aw�������w�f�q���:|��\��?��Q
��J���=0�(���w+�K���A;�5.{~�=%��( �n����Ck�#��rFw��M�2��'|e�V��.���U���[�?u'�Blf�!�fA:��Aj�ή����t�� a�� ���*@
%Aߔa��q��qY8¨T��Ϻ+wZ�Z��Rz�vZ���x��(�\��A�\}4g?��}��o�}�j&�S�5�l⫇#��`>[6����c�r�5	Lp/A�w �&F�,0ɢ��;�<R�`�~�v�R:�*:�?��0^?���g�J�oe�� &�ֺ�N��qC����B9
��i�rEd�ɔd"�����J=ڜ�Vp*
��B�H���0]�X�F�sp7 �(���L��~t��W�K{v�xAY)�壱���!��;�u�Ou۱#,=I���I��&�v�,�5\@�$�@�_%� f��Dco��d[P2�b��|�ᙡ�0C\ ���"�,��ƴ@�򈓉���b�x`]��'x�H�7�C;b�-�6m����:ӑZ�q���Q���0���|�:�
�?��ʵ~I8@�~��!h�@q�^�\S�,�	�Nf�c�X�
^����σ�� �mЖ$e���x�y�]aD׵��?�������Hm�v9�w=�mX*��e��Lj�&�軻�h�1teD	�z7��$���{�-��k/��v+�c���]��
��u���U�W����_��O���.2�n[�SC����ݿ~C��-y����'E�3�, (v�c��P���/��5\��B N��Ї��潡�� ;T��+�?O�[� ��J� �H"�B��٫�0���_�竫b�Ӏ�>����[o��;)�鵯\r��pe�T�Z�|�6������\)f��;��:�1_��ڊ�ɝ&��d�S����҇����c�d��z�kL]8�M|��o���w
�/Gʯ�G�9?A�L���`X@���/�>gi#��Hf%�O_�eI���SEhDj'�B`vB�K��:�
gM:�
GPt��"��|!T�7��k݋O�&9v-�X�m�T���}�pp�O�"��C��	$�(!焂��<-� �?I-�e*t,F����(���<o�k�� �.�̀�}_~��r��\KjR� ���pXf���4�I��-p4#,p��dS�}Z� /H0��^�2�L��tJ-X���I�U 	��]�/����0"8��0�3������Nh�i�y�k�ؕ�g����ͣ��ϫ`��-�M���"k�\��jo�]����!�6�=�5gf��</�r���*A��������d��%����<Y6�E�$�/g�=
/XS�2t�00�+/��&�����F:_@�0=)i�GN��Lʼ��`�g��\�1��|�C�(͈nO�O�L�>!�	���N62�`�׷犗�@1D�Ot"�ȑf0-2��5c��"���;U)O�U�+���V(÷�)�nT���r����������|�8'ţ �#��\l<r�WW`2���-�9�����G�;��F��0��p�>����e��e���FT��R|�����:�	�V�!�T��_(N0�;�l��o��c/f�9�F����!�&�������d�Z�z0�.L�--���������F�M2���F5�?9H�t�<j%��XOT�Bsw_*ʩ;}�f��&]��ѯ��}"�[���h����)�)�j�Ȋe��U�1n�W���;���0~'5����uN߼}�ȳ
"�����mը�zgA�AS&^ ,�F��������n�+��u�PK��*"|��G����X�i��%��j���y����[�c����0p�jC���-�[���K󘪎6@��Q�,��Ɔ)Ŵ#��ꞡ�ٸQg�󝧣08�¹6E4ܕ����O�m�#d(RD�z]/��^�ox���n0���]+R��ε����lr1D#ݜ�j�x�ʺp=��)�8g��`=Mi}�p\��4|�?��!�5�I8w�	���� �-5R���]�pRP~�U�O���;8�m��~����pޙ�u`��9
t����~Bܗ�Z��w�;}uu�D����k�^(5�Uux9}�'٩I�qA�X�	��>N����ug�)y�D�������O%@,���K¹��
��\��ݟ�x���L�E���@XI*ͨ�Ճ�k1�����:�Ls�,�_��?�Y�%fwY���D�CUE���	�ɔ7�?=O�Q���U�a
��@���Enu�އ�:y}ԥ�\��c�Rh��"���/��3���Wz�Jٳ
l�f"z��F�O�0�c:�=m�I}j�XM5΄�-
��Ϟ�[W($M�Z���n��*1���o�Թډ�&]A��p�iĕn��%��l4��X�5!�!U�e�nj�T��OMT��9M�I�aRa���Y�o�@x�W$�	F�c,��3��H�k2��+o�:�