XlxV64EB    15c4     850�6ghS؂�O�+�	�#{��@�}��=W9?�������f�y�~:�)��_���qr��iw.�!�}ʇ�>�3�r3<UB��]7�OKq��]mR�����jx6��.U��|����)1� 7v\�,BsQg^���zΐis딏׮��ހ#[g�Ű�qғ��n�Խ�,���c�B]���G�kR�1%�D+X�Y���}o��3g�m�%S�cI>�ۣx�gU���+�4y1��2Ɩ�S�Ju�����%_�����`���wo�� ���{p�9�ihL :�i%��b8ޘ�;W��Q��1~A�Ē��oƎ������u>�~|�a�u��(�6�wL��̫�_X���Wf�g�Y�x*�N�t�t�ZY:��P5�ZsA^��L?����]=q��t�vR��MjhD�����#�<�<���θW{��Օ�[Q��0�H� W�9j���� �uKs�	V ���7)dΪ���qD��.Ȱ?y����	�4D�;�"$<���K��*#�!��-�}���^�\�ij!N�.�o '��'5g�W��_�Շ���?{��_[vIG6�!b��@�y	0��{�~�m��p�x
�;�r|�$7#� � �+�A�|<!��B��̮�	��K�����������ξ����҄�1�E{1�e�N�Щ='�w�p��
%�|?���7�ʄ��'�  Y��o�CO�#���(��N͖�	6����͆�|Βaٴ�����o߃2+ph0:� #�[ěgJ�P.(Ǘ���'�C����c5̐�G�>����,���������″�3�Z�C�<�Y`���>K���m*$Z��|� ��.8.�Q��n�Q d�?������li8�#h������8�,b�[Wc��o���HFJ��>��B�G~0i&,����� ��[�zнz<���3��`>��I*O���o���c7^�x��(�'��:p�N�>J�'���u�+0sN����C���)ޏq�"�<�f�jmi�����-��
�����)��;��)�dK��y��>���a�
��O\2��#çJV�N�6�ov0��09��iߛ�|�����huw�-<� -�����ѹ�&�Õ \{�����Gw;�Hm�Y=��X�����7�yϧ^]�Λy������td�0JMπ��l>������׈��+�7���2x%�����N�y���7�j%s_}B��� ���:?�+>l��4E�r9Ū��bA��۴��hU,U��#1�*�� X�^�D�9�ƥ�B<�(:4�K0]`:5,����z����vݒ�1�u���-��4�� ��?����lQc�e.9�����?K�u&K�EC���.j����Wb�-~�F��d�hJ)U��r�k��JQ�����P�1EC��l��� ��f�+|k�&.�u;,�:�9wa����`Y��̗��
����}W�!��|�׫]�o��z��r�S�~�}R�����J�\��|��"Е_��[�ś���=����F1ٖ5#.[9?q�$���;��Ih(��� 6e���'�9��S.�S���dB�9ve���~^8.&}|�MEV!WԒB��oߵcS�d���g�����ꦌ�~�ٛ�i��Y�����Q���q�7N��c�����9Xu�r��4�<�=(1w����a���*��
]a��k$%7��~�x:��>��	���l����skk-�M�f L�d�(���^A�`jg�DI��]<xa�N����B����~y�R�V�̜m	s9��� ��\A�)�e:=���G4!�9'}h�e��/�*�h��K¦Pg>}$7r�3�rx(��JV�=��F�9��K�3��dɍ��g���D4~h����1�y��;��̒2ԖW�o����B��M��%i��Ō��}=�8��%�%�Ӈ ���M����ډ��aJ���;�s���@���@ԋs E����C��q�o�ךg1�O��LR>&���Nc��@J$�W
RJ�Q��m*����<>�!4����$��o2IX9}'�B�u
h����y��h�`��