XlxV64EB    2395     bd0Wr*����y\�S��Ȝ�N���>�鐈s���֥'֠�޸��cO�R|l=5Z��J�k�9�<C��_�n�a��_)!�Hxk�$�)���*t= � ge�ԡ�l��2\Z�/�*����?φ�4�p��D������>V$kI�A��(>@h ��a�^�g���zv_���l�ܩcԆ�{^�m����?q_M��t��5n��b�m���g�}D��SH�.����b�Y�LY�-Tm
h3��� r;�hcC��)3d9��y�5{��ǼBllNܿG��Ɖ֫�@VM+�X��B��V ��h�7���0�=� T��f�N�ld��:�*��Z��1T�"ƥ�	2���@�k��K��g�ޅ@�����������\�$����B�4!T{�=��{�ū��O֭��5����'������9N��5����^�yLGRa`�����H�����m���u��
���=�8	���"�i�
e���vL�:��r��PmY�JΊ�>\����xKHmА�v��(�(4-\,#��ٯ�/�1;��,YxP+d����?r�m.���O�T���l�(p�>�B{o߳Qh�si�X�ܘ�*@���d��.4sn�{ߩ)WԔT�׶���P)H�3m�|&���7��9�����N��9�������V��S�7���<�E���K���Yd&GtƋ�1E��Cya��"B��.�i��������e��6\K������:����QP�_Ӄ��j���ѝ�iBGz�J��K-J5������I���DAfv�����_̈́��t�>��O��m����ڡ�-}^Ր8��zq
7Ῐ��%2v��$��NH�v�^�Ֆ ��\��"�x��63��d��!y���L���$�����^p�WB�(�Tuiaf��^ �.�Or�&Im��,,%!nX:����/	_R��)�M�'��2�eg�QѢ�C�e��Ǆ��=�s!�/��9�i�*8g�^�j#NshC�z� �t"��if�Ӫ�a9�d��8RX��d�})?�����`o�x��^��J\B�;�>X�>`�^x��<g$N�0�}.���ڵ��#o�h���Y�e�̎N-$����tu���cSl��ʮ�;�)G��j%��س~�l�+@��Y�>߶�b�k�@������0����e�#��i�.�:8��HxAG��U�<�=����2d5��'�	F�FFw��X���	���DTk�5�7nygu%�� ���J"�PEd�\�	
v��	"1������z�,N}��qΜ��f��jL���=�&�Ê�}��<�K�J��M�h��S�̢�ϓ�*�)����+.[S�AdIE��t\nj=SۡR�JK���xH�ٿ;itl����O�zD��I\���^O�S#��(M4�r&�v�JP���@�9�V:�`%b�,I��Q�MEz��_t,qhK�g��p��%Z���B�'�&�X�;�f��Ȫ���K/����@e��)7XV�!�� �'zS��j㴨ޛ>�����R��� �j�}��*���o��*�\�yb�#DQ .����b}ٷ
�����ܢ�H����kM�+��%�3	(L�o�� Ɯ�g"E����〻��;��"\�J��,�b�/ͭ�~��t7�M,��6Je�HcEx<��r��c�͉M��Ei&�N#'�D�y�{��O<�<k��<�/�o����Yq3�Kq�A3F�,d�Z���p? >��=�Z��3�?#� ��EH��`��{W�IV»d�Q��g��4_nn����`]~oF��=ϩ���E��4���^�]��+�	e|FiG�Pzd���?��Ȕ�=�e�A̙2�P6,3����G�ű̯����,�kKZ){�֬�&���h��=2��/i¢T�N���(+�����$L��**�nBx2�]��T��)�I"�����I�@r%h�jI�ܰ��V{�J�h�g5�i��ԷͶؼ�'Il���\��y(-�����u'��X���F��I��[$�ܿ��BP�[>�� �cZ3���_A����A��>�$�O�2����"���d�QXܒC����l6������6s7y�������{4�~π�)�2�M��88��L��8�V{[aZ�˄���Q��g]�4��{�>v
��Î?�q�<��Q�	<L�P
�S�]y�,�M�A >��U��f}1�֥�=sZ'�(��/��\��?J�>e!��:	?FY��~7y�������:a)�x�����_��|ð�ڢ�|#�'��@��.7��]z�]sO53R�6��-5(�������v�gwޡ�\�N��+I���(�"?Be��U��T|����ծ��\q�_$�2aQ����6����'Ķ������v����y�i	�?����'KP}��l�v~,$�42X���A�J��M${�֕�/ m��ɘ�#��0)�I�.�Dr��Ҙr ��Ҥ@��i�ɷ�9ذ���-~Y�S��O_'�(n��屮���Xw�Tƥ�XK�ܖ���6;_�!,+�a��@�"���;b^���K-"�CMY��GB�=3�?z��:3���;ro:3����L�|T���*��NFp�0]�:Fz e�(����P�b0���j�MҒ�-�PQ��q�ˊf���=j��c<�W�6�H���:�.�{%(>�)1g37�w��X��yb��)����W{GF;�:��6�u3	��:�P�̂n�v�Ny"��[?,^�T� �����ʢ (T�>!E�~�^sT'J�Mp
�D�+�e�R��,���b|�(v�Q��f�<B���[X�C���h���;q��/�j0-!Z��#?�80�I��("Q�i� s��k�g9;y���򌧍J�ڢ=`����d�"�۬�,�{��3
�� -�8��c(�9�Uh�Pg�~�H�