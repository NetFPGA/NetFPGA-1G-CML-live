XlxV64EB    2c41     cc0��.F������1J2M3W���="�t�R�D=_�g�6��z���7�H~/xaH҂@Oa7N{�T�p�b���6l�CMf�y�����m>Z�/� ��4�S�`Qݽ	gDOX1/��v���H�4��O�<R	-�*�c����[Y{���T|��mU\Z?��!\3��N��[=��8om���<	v�O��$V�(icЬ�!?� �ڎ�~X*�V�*h�����dY!�9-f�Ӵ>���K�ހ.���#��E��_������"`�7�1������R��8������R�GR� �ǢtF~�G�R����s�~#
�M3��m7�5����-����ξF� ���]���Ґ�����8�tv͘h0��>-\���.@.Ҡ��~̌*|MHѼ62	 �Q�Gc1�Ҥr��ǓVUM�¨$A/�Yp���>�-XWKa�^5�bE�+�Wj^̠�J����ۘ����R6��J�Y��RxY~�0������R����8�i�qd�/�L���;>ѝlw�\��s~GW4����:�7��`pk���R�9�$�AxMk�q���9h�ſ��⶜e��G�?��>c�����;n>��a���cܫ�Jrn�!�N�5<�}Z�Z�����5K���pB]��0�M+�Y����n��ת�o�9t����� �p!p�~�c���.�����-qˇ���x՛P��B�m&BH��r����m�r(��v���R�ͽƢi���yc���U� _��ZwW5�QV���k��ׇ[x�9	�܆��@P�>��+@d���K����˘M������F���6`#wJ�R2_R���M�i'��5j�*��(�4;Bq� �iuX�����}�Y����N^K�@�xq{cy���<�ϝ!��	n��8q`��1���DT���
4c@��f�c�;�R%�qf[�%��ԱU%<abk�����x[��f�vQKE�Z�n�2|�~{Jc>i�~')��\�g$���cn��)(,��T�q�O��>��0�ҕҺ��'0$�x2�=�?��L&;m��/-�lhK�C��<��=�S��7}efF���#�Q�d�_�'Í���/g�j��&D��0��*E�+��Z����k��-� �ѹe�p<g4F��bYK$��C�(B��+ aZ��S�nG�������k�cD���c�4�B����C?4ZOOP[��ju�[���@  ,�Y��=�p/mH��s�"����S�qM}<m�IG6�]��!�E�0b�:35����x5�`a� ��C�P��x{�u�#d�G}�.��������������AN����>ۑ=�{t`�-�q�vBڃ79΋�����p1J��T �`E3�Q�T�fd��/�2E����G"��5opf�=�$gC�N�H��U�ݼB��Z+5QY鯥�(S9�g�z�����U/�5���<:Ga�#o�Ϡ���,Ӓ<�nЙ��W�q���xO�t�]k���˺��Ww~TjY֢��[�*�i�M����=-~��Y�jy
W�X�A��!>�,x)Զ!f���z7����Y��yHMp9
���A/�<��N�H�k�Gݏ��
����;�άy�_�~<+j���i槐לd*�g8&i��1ɇ�+uD1$�����$�aoL�q�~�+�T��k��[\ �@���6�ۖ��/����� C�J� 9r�)X,NیѺWAӮ��sAON�)�+1��[{�т��k�kz�]�����d	b�c�4!�	�t{���>��������ZM�y5�6\U�9�b�'��L��{@��Z�A2��0	[wCĉ�[J�|��?Y��a�y( �]��m�t�X#�i�^�~CZ�֐(,:�<fV�	pD,i�W���F��%��N�L��?���W�Γ�!�I����G d?7��X%*G�O��|��''�Z]Z8=YQ[���G�bEF��ϸm��VnL�,wb!YԞ�D�[#�X��o��z�^*����>>����[ǵX92���Ţs��U��e|�����/�q5g@\������S>��k[���oO��{�MR���k�5�Ƃ�!���>����/7�y�<�t�?b� �|K��(��~|��9�5��~>+��`�Q�}��dIUA�G9a�����D�@a��fL��$8+ ��l�y�sɮ��]lx��pxj�`B%-��+sq�g��N	}�ػ���r��9�r�d�[����2<{��/��LIR�tf�9h҃��y�L��#��
0����!xio�b.s�&ITf-�mҷ���r�F�!%ǯ�LGhb��R��
�Y��U�F�Ëx��]�'#���w�l=���,}�~w46�U }�[�.�*�Q��C�$��g�E~��n!��Lo�i2��92�g��h������yi����y�E[������w4�j���3���}��M��|{}vj��ӄ�x"�h�״C�������W�	x�t��mm��c�K�Y|sG�VZ�����9 �g~^z0����~M���˒ ����	���l�ϗ^��S�k2����B�'Q�{�A����&^�7�I^4�o�(l�);o��p�)y�� 8�nM�����>e|��K���b#��Y�r{�Hu�5n��1ݲ~�+K$%�H.-G��t2K�[L�'�҂P�}�|��w�W<�1�D��a:� D�� I�>���<:׹��:,��{���CF�גZ�ZM2}A�0O��l������p��4���J�2$�E"Zf�� զ���tz����%{�����ũ�ګ����E�e�"���e��W��m��9=�Z�W��V34jb���� �Є��c���ٍH��7B�ʑ�ށ��߮��B^_Q��o�#0}_U�l�U�u�<�O&��)+�T��Wu7&:��MP-Mq�-b�9}
������h��V\����Pq��^�.�Ym��xA��?��HYcw	����~�����g�{�ų����꿵W���w��t;��LJ�j��.�{G� �t�㧸��j�z�f[��V�@���#��ɼg`�����6�J��.9���8��`�/���m��=vP��T��M|�e ��!(If��)�t�Ov�m!�?����G���n�+�b��� ���Ƴ9F.&=;S�V��cňm�ӄ:�U��&w�aM�i���7��@HY��q�w���m���N�7����y��0�"ʤ��

��eQ