XlxV64EB    3ef8     ec0`������;ti�/�AB����K�23�f37�*T`�	���FD�+Jg �_�Ĉ����.�AG3�fZ���g���
��;<� ��~>�2.��>g�Oo�*b�:�U�C���E�=�C�f�WD~����XC��>�w ���7kٛ��D�mǓ=c�(����5:��i�i�	��f�&��Q�ZvU���4f:{���Cn�0 ��з�=-��	��8��!�9����C�g-�E�:}�6�T�-* ��ubH�� $WQG�[����������J��D/��)&l�(j_�����d��B�������wn���\��)�~d��+�/�dv^fC�{)��P�UFea�9�@X��F��Ck��
�}x~����%#�Fb,�Xv.\~��g[�"]�
�@�ܛ�F��ȭ�a 8��W:���9ű�O&��Q�����H�<v!G[_5���T'�rTt����q��j39��./��0|��,���%@s�[U��z�Ga�*� ;��#G���(�&��|��q�/�{��6J�ɲ�F3����)�)�ՇQ ��$ta�k�}�޻F�(��֋V�B������9���L-�F�Ze%���a��V�Wd����<ٚU?`ׁ�~�����c��2��.%p�7q��`8X����]}�o�q@,d��d6.T�0���H���8���Bu��q����,"�����k�^\6��VX�멷%�~��w�Kr:o9��e\��N�/�No����ξ�Tu���i�.���\�K
�s����	/D�@�}����@���X��ı���3H��[$
�/G��ִdK�p_��|`
�[�CeR���1�y���/ȵ��V�[�bnY/�BY������&΅�A�ў�J���i_F�1����Zc5��]�/���߳~h0�K����0ןAe���Q����Lb���T�=�H���Y+nN�ť���q�ZL!H8_�j�1�����=P���i�yU"Fݸü��@H|��d�����&I�Y��֒3�>��w�j$���ܜ����Bn���Ϯ�vu����%(�A� V?�`Z?����V�?��!�(h@��uhZ�orx@n��u�@@ost�ʫrՍ�D��U��.]mƊj´k��J���2�����.r:?��Tv�GPpO�w����_[�Ɍ����Ss���kR����[��{Ɖ1�Qp���s
,h�*�{/%�����:�3}4�,���{�}�ቑ��`�m�N "	�� �{�h »`��J��Jw0��w7�Տ�p��x�b���~�|��j��kR���]*�'o���v���l�I�#Tl0˙��*ﶔm�u4��I�L9f�e�{%�F	��R���[���'����e�
ոB���r��;S�IFv8�|����>�*�����ˬ��Bl�!�C�γ`sv�)�wG��<�5��׶z�G�9X��,cū��A}2�K��ZA��a�6g�����gRXP���#�&�t��Zֽl<��a�+y��0i[�IL�@����D�k� ��P�ܻ��@�v.-�d��e�Q��a �l���*ɑޤ���4�o,1�)��cɠ�xʕ�T�ۨ�#m�Xm�W@���^Oe��e69Ν9(h3	��++#����;�X����*���p+�ы�ݪak��13%v���3�w��p�I�=ծ>�v&�l�<ʆ(��z�|Sw��rNwr�lH��)�\ ��^�(K��D�=7YB�dA�o7�|qg��|8���p�RkB9�K�$�����&T3����H�i�y��!�*u��li'@�H�C@.�㈇��xV���V�s��LT�o��@#1W�b���vf|���k&��>��	xA��ʳ�)��Nm\�+2Ȕ��X����ϛ�$�nTD~���NK������=�znn��*r��`\��g�6�&�!ܒ[z���ѧ{.`X9����gW���B1�u��i�p���v�h�t�!�t���
#���7ȻԦPE��c#��ӰNz�ȅ���|Y� ��53�+�����F�.�[�D�X�/v���@���̳��ppj%��#q.�L��M��<ع���i���n�f���^����׉KȌG�
��T�i֥+�
c�� � ��@dKI����c�:ϱ�-�3����#5���&�m��<�|T�;����_���࿁�C��JP��)IZ��G�iO�?�@�H�1a�%)���9;�?��b�|R�3C{?^��B�z�^��	��z�d�f6M�%�+&�T��[�r�(�Hu�7�wC��qxI��!� �Z��ت\�{A�� �m^K�=v��.��<b��+w��@�E6E?ݹ�A0�T�E᳥IK�৮j��ß�Z�5��ª#��!C d�hB?���dp�[��O8�;�<��3�ጤ��k��-�K ��y�d�7��X���L�S�R�Z�ld"�=��ݪ�`]
��Պw���E���VؓcO��"9j�:8-c��dP�X�g`_�5b6���~��!�fiR��6
R9�FYW����JGA��c���p�Q��2$�@���_*w��\zK���{J�81&��9F�w'��o��$����\X������ q�àD��E[$��dKe����y��m�R _�y���>�R{��[4?��#�Ȯ=W�xB3��Ob
��������������ĩqc=�C��Ҫ4�n��_�����|�S3��<��ԕ7A�U˳���Rw]oV������5)v�p����[�v�:cP@�h��[w^EK/_�غN��XuEF�_v������^_�x����C�#�2�d�'0K$�{�xIV�߶���ࡈbF�~����tg������hs��2��n-��N�ͅ��u�5_tݑ��j蓺�Ȗ�_œTK!!Áb=�/4��5�_�ky㦠�8-O>FWp��>������[�<�j��9=���7�o8�%Μ�^n�y�px,9��׉ɵ7�#i�>i(Wچtj��qT�a��f��Xz����46��p�t�%q�3l���G�����/#�{�e��ٺ���zW�ݞ�g?���l.p�`���R������,����eO�����\��$���ײ�T:[r��U��%��K^Z�B)Vl���d.�>�q�c[	��&��$.��p�˫폆R�x´���@s����s�#�7�6WS+㍁];�u^��{�������T����!�T�-I���
c�̖��G�z�	B֊���2�B���(�Sf�ը�6m���w�����fi� B�]�Br'��S�N��}���hC;ay�h�b	{�g���� ���M�d@iத|\�eg��>J+���1�O�7Xd��U>��!j_����G(���\���{��T�@�~mm�ז��Y�R'�$W,?������3å���1�����A�j��h��l��z�7���� G�l7��w�L��tu$�*�t��`PL�Ӯ�+eiՅ�@���Y�[_7&%I����/�ԗm�HB����,8rk;��:����%^�������G�1G;ZZUk�h�qZ��Ԥ��O*�(͵pj���'��Q��Z$���{����P��d���,ɟa�I+��V�%���:�w�LH,�xM��`x�2�$/�