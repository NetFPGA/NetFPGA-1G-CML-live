XlxV64EB    88f0    1f00saf9����	���������b�[ĞH��J�0ո��	�֨��Y�X��:95�jJ�0�(���ZA-AU����x����������'-S'�i,��8F��?NY�nx�����<�$t(H����E�a�]���b�N�8˓l�^���I�K� �la�<��h ;� �4	yQ��QS���Bܣ��C�����Gv�W���o���c>�6H�IQ�W�P�����yF-m��uȧ2[:&0 V7]�AK�q���!�:S�����'�j"E���r8m2�r�����A �eE�'w��V��$&�r�g��З"1nu�y���#�$��B=]���6�F�� +r{�e;���Z�V;Y񳢴I1���\�kD�~8y\��\n��w��-A)��n�i���3XU��T��d��ֲ��蹓#�SV�!1@F�����djl�ן���E�C{��֙!�� ��3�!�?�D��2Igt��(d�0SY�/8�KOC8��_��7W���@�ڲ�<���LOqʧ�
P"$5�#���i�w��{����c���m[���A�W�.�3<:��_�����r�yØˡ%m��&j��a�]���W1���A~ i�/�S��I��@�zS��߯��C� z��'T�?��p�Sa���M������_[i�xU�3(�ImT�1�?v����.�������������a3���8r��ُ��������j���F��T&�x�<���� i����W�R�u��q���p:A�����b��S�[�t�ڲ�ID���P�/W��2z���z��3,�*@L+���E��,b�u�� &j�7�d$�c�7� a~��
��g��%��P����d�����X��4m�j}�Q�P,�ʓ�c��;pw�����R����M��^A�«��$���V�0�9?f�-�����T�g�L���Kۑ�p�v�>c@�$J��QU��*/+Y��8JCu�2Hq~���i^6��O��;/��+.�ǲ+�;�kat�y�r�������l��c�EnPT�w�f*�5�K8��K;Рa���7zt���t��w�^V.�%5�"����7����%WąB��}/����s��X�{�*���'������廅�/��c�hv�!���k]�����[��΂S�Қ���0�̧�)�:���Wߟ�f�M�at�όd����ہ��|�7�):f�������b�>y��BXN�9Z�x��~���ni���_�)��ZŃ��Š���r2z�t5EPd�}��:�~�࣊�\����8l��&�0�X(�g��ҵ#�:�z#�Vs��u��dΆ��T]"[��Zֿ��#'\5�>r�P�q��ap��]45�ck�)�����В�N�!FE����~��rٹ�補�p8����{,mǔ�J��9}ay��`
���N�@Ϥ5I@�/���>���!~����Q~pע��4eBIK��Vn���N?ےn�B����f���Cx��\{Y$��S�:6��jݕ��!�*�pA�-;�cQ�� �o3�n#OoV̻$/k�a'��l���pl[3|��n��~�a�	$W�I�7s�m$*7dѯ(�0�&G1�l�u	1���ڏdw�8��֣:�����"�8{�,��^��+�ӭK�\M=R�����! �E]X0a�Rx,GM%����\>�z��!�C�2iTW�Z�����"�Q��S��ĺ��AA��ᇭ�,L��}_�h �������U〞����A�5�L�~�5���T�p�'�V���tt��(�g[������Ვc�"�H�rP1�e䂾���m����FQ��P������(�
ﵻ�vx8�a�y�Zʖw�<<]��у���V۝Q#��nQns�J;^L���Re�O	��v��?��?;M_T`�x�Yˇ���9Mw�ޛ1�Al�T��N�+�J3��u8&� ���Fg�̆Og�=�%�����e���;��hv����v,/_4�ԕ�-�4 �1ͼ˿(G�{�vS��1_�Q�a=E�.h`�� 1}��nc����0?����AzI,�EJ8p��>�ڴ�(2v�x��]A�t�x�y\G������R�^�~�v��S��ٛn�"�϶�v6"���*��R�xe�[
L2)��,��0����G���P�+�Q�tB~,���s�Ӑ�Xҥ��Z �ۢ��[K�h��-A,����1m締@C|3��(��L�)�}�I�7Ө�X
�aGЁڔn���"xi��Y���h�Z���o��D_��f��Hh��9�
�B?�}'�&��I�]��������?=\Y��W���"���}T�Pظ��.5��i�(V��<pH��/����Qh�܅�^3��y�+�Y�/!,���]���`�����Q��(�QI�G��9��զ��^�R�,���BU���M��ȷi>�p,�-��eI~�3x��W��`�я���==����C���Ƣtb$}����)��d?SW$�hAJ��?�`H%�	4��"3�V{0��_!o�r�[�OA�5�$H�.9�������g���02���O�-�CM�}$�YR��^j��9>"���K��f��|� ��'�/4��m�;��f�`�u�2���=6���F�r�2��}���[���(m��`T���َ�kHDhGX�X�Rj+���n�0�_	�.JA����^?����W��V�nٳHR�O��m`QA��Y6�[�{����)�a� �y�銫և��ka��/F�L�S^xV��:�<?���w���y8�	_����xړg��*8ʢ��˜)�j	�3O��?K~ٴ����8ڈ�|�w�Iz;ԟ���锜�ٱR ��7�{B�^�i��ƅP3�FE�f��ܚ�LD��6X�
�*?TW,�T�[��U!� �ī��C �M�_��=��b����!��ŧ�y�{��LPd�@&����s(=�4O�l�A�@#ᵯ�h�}�C�uE����&��i��j+9(�tګ�ƋP��!u�fq�_%hX<�ɥa�ы79{h1=��M)b:\B=agx�(�5�y�����Ԁ�L^P�2s"X��iu@�ޝ]EP}Ä������±�)J����>$h�B G�G��C2ٸnh [;�4�M�5��V�Os����y�Ɯ-�����@2z����	����g	 �a�*� �}\QإyIt����S���� ��g���k���
^cX)���I1೑���bp��?�wsT�R2[)t�����u�NH�uxZEb^;>�{j[Ώ�d��ȗ�U�GL�TLH�<��B�5�������`�=�n����pӓx}oj����P�WD�S%�|7`3{��a�L�:�骮���A��U�2ˢL�_��<�˲
/�Du�fh���5�Y�&�{&�*�]?�uX�?�ly"�u+���iI��#�	�E��U�L�('����8�*
�s��C��V�~6h9���z�g{0OKDf�ٷ��D�m���u�0��4�ɴ���xL�	���ep�U�=���U�w�{���2�H��I�o��mKË(!�����ZU�����"��ܰۚ�VŪ�J8y���TA�x����[!�qx'�tEeɦ��'��K�O��m��$���kra +>�p��q�]��V{G���3��R�7�yM�B�/�~%�,�r:a6����Դ~4��5m?R�Ar��h��
M���D���������s��v#v��x+��in��
#��1��r�g�'�tZC:E�'�`^��y�B!H#�P6q�@1���r���_4<�1����s��������j�1�l���"�M��n���Y��d�2jB���Aos;�_��?�q�љL3y C�`�BLs~j�K<�E=� zH���$����?�n�f���[=0/���c��a����n�RIe))��xWr�
�����y�%Jt֋p�a�W����۾@3%
]H��{gm1�����)z?�pJRA3�([u�;}�� ���2eo\#1���*3A�	j��	,� �9ڊ$�|�E���8nC������F�~�?�V+e+�*�H���J��Q�׋�Es곸:� _�{Ek�|A`~�RZ༂�7�f��%1�(`��9�����X����QB%�*��⧰JD65E4�����dZ�V�mHb[T�������\���h.Y���AɊ#��+ي������B�9$h�u����J�
 p����k��O�Q��o+:���hۜ��8��{�GfY>�tYK�����8z����K���Hi�N&h�i�zX��&����@��J�
� ט�u��#�kC������R��!�o�\n�Yz}嬩�Jң�_�(��=9qXt��<�$OS���̽2��jz:U
�_�T^S�T	��RnO��'BLy8�*7��'��oO��R�O|Y�'߀����C��dJ�{�?  �қ�yR�s��	��]�J߶��$�N(G�*���]�V*��W{lA+ت��L�*:����	�3�"mCz�(2c����۔A0	��p�Z����q�{Xch0	H��	�Kp������*ݵ(G�T7B2y=u��e�IqG�r�<��sX$�YB�,���\@ef�HN��t���ҫ�x`6Me�lÙ��Gy�	�@����uS坔Z2�Τ�]�u�'�R���u������r[�ܱ�c���V#��S���2��2A��
������} �{��Gi���y��$%���\p�ȓ�aZ��)S륖�T($�t�kͷ�髨u@�.�a4�k���A��f�1^��M����p���f%��U��9��f���̨rvP����	k:���Α����a�p�Q��[l�oZ����35oJSu��������' A'�0�mkMΥV;���'=6D�
��R��dc�?�@}pn�x�E�I�=�6d�����Gcm]u�|-���	�l �Vtd�u<�d���{��
��ѧ��F��3�3�5�r�9�eV2��yCx� 0(5*ޡL^K.�y[s-�}�3Ø���⁔���>YQ��
��_5	`�Ø:c��A���n��=��@�:;E��#��R�]�ٚǮ{�]���H��E��@�7N��V�]��C���c��jf+FN���픵�n��n�B�����:��Ш�@����^Վ�)��YA,����d�C4��t�=���{�O�8���~!H8>���lx��R�ͨ�Kp�_�
���?R�Q0�p&����$ ɦ=�gf6 `cR!�����\��g~�`V�j&U�0�<֕�-���?g�s��~M���gк�i�R������XFm�T�D�ݥ
�$r���T4��uEc��=W�����p���a�k|F�HFL/�򸉓���w:���5���P�4�_߂
��<��#Ö����Ř��Y���՗��j��3�2W�4������Ք{ϵ���2���D� 3���
b���fT���Ac�<�ɩ�L��v���UN<WB���$闷	��U/����h�CBss��yٷپ-Uq��lM�c6QY񶄙���=e���G����٧#�犵���`��*���_�Q�Ʃ	�����t�H��{�T��i�q��Qf�x`Jx�n�QG���p��>YnR��c�����U&1�a'B��-�O��Q]�:��=��&C�<� q�-D�F����9��,���?.e��P�w�;¹,��P.��f�LYZ�9f�ǐz��:���~%0�!����f�n駜A�5��e���_H1Y�.�!���}.��C�a���+3�5��C�� -��� ̓_g[z��v\�I�&�C�pbx�V����^YF2[����>����31�ىc�1:�������t��i-����J�"��1w!���,�(eV�/�{l������i��:�l�������?��o&���u@���[ms���T��8�~�x�7y�[��0�?�Ý��o�ؼ�`/y������9]����v�Ht�''��X�)pw`�!�H��v|,��Z!��O�#�Ұ9�u��iѩ����VCV�Yl �5Xr�]�`�E�S���r��ڕ���:�0�J_��9�x���g� �3���`�i`��q*遰s�����H��Pp+;ݱb��_�_��2'�t��O�0\�~g�ë:x{�-lC	����B������v<���_��땃B�cYZ-ܷB耬�e��Spr�f�rS��ʱv�N��&����z�sR���8�74Bo����^*�}eI»w ���<�Y`�*7w\���X/������,N��RFn����0�WS4;����;��'�j�l��Ks�)�S����&�A�k�v��9��6�B���s�i�⯳��s[p�+�:�����L�iܪЌ�aOw,8�`Kx��3j�;�c9m�Bj�.]�8��~_� Se^ �|��\�1�&Eru�o�p�#Az����z�8KQ�S#�4��l��0]������0����q�ZLi!}
��L��/�Qg��%��|����w�18P�\S7�4��v�Q)� �/CX	B��vg���]GN�-��@��-tԆ�?33�h6w�;�E�����~p�q�e�U+�Q�cm��~{�E��=��f���y���>����e�q<������a�.�t��
�t�_��
H1ԡ,������sg0��Y��^c�K�S ���aw@���l�JJ��o�QHCo�KA�Ԅ�N/x����Ě'�8�_:
!�#�^�����L�ч�y����@��ua�L�^Ř�D`1=u<�tI�V�WY�
�9��k�]
�|k4%2�mp� 
/���̍�l��H�~B ��c����YB6u��zU�2��QUF���p�1:��+C=��p�RԂ�d�x[�i��<PY�KՀ��g3Ã�	P��>�
���'H�X\4���ݬh_>�4iJe/&�z�V�iv��d�*h�+�C���nto0����FIm��8Eu�O[��n�6�{����U<t��.m;|!\q�=�#
���u:�6��LA�YM�j���8�:�!����0e,Us�YJ���K�'���g���̔1�$�r���4&��I���b�%:�Kn HږHyJ�{�V�ӆ�>���@�+����m?9�D����8c��`g�݀��`��&Vl���g��X����F@����X5kP��O��o�8���gM���>�fd�;Z\S����jå�+���,	�N
�ͨY*�\���7Қtn���p͔o5ͬ^�8�w�Kjw�BTKozb��+Z���_̧��/�{~�W���0k/���d��DyZ����_u��Ź ��.1	����WT�7	,�JHӹ��w�V�Q�^�ƕ��۫n��w��ˋ.�_V��~)E8ErF�D��d�h�s��b�1�|�#��8�BZ�2���\����E�l
L}�+����\���7T��]Fn�f�r�2��L��f�W��j}o�A���s("YB�]S*>7��2~�|+�o��n5�<����z�Ė ^Э��3���3�^ʴ�[%�ek�ف''�cn�3J4%��(W��Bk��/[��~�ʵ��ܦ�IE	-Г����8���@�\���1�5�V<���p�HD�gu��mz}k��8=�Bt=S�Z��m# 	,�[F�����DK�4}┧�v`.T*Z���m=Y+�S��O��kT�)a��B��1b!�^JLb2�,�4