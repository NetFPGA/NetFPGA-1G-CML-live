XlxV64EB    2a88     cf0X�����.��Wq
�ūy�F�G�-3E�<5K�]�+n��2��s�RS�ɉ�׵f��Cg�X��Ï��Z�L��0"o�|��.�i�O����fB�^72C�{�h�\y|r���8������1e�'�Ѭȇ��E�s��#�޳���<��0�ִ�19Q(	���X�F���(�˸R7<��#�b�O��/p}1�&bx?_T�	8�1�۷"+����r�����h�Mv��>B��v�Kl�o��C7�H'�q��U�;(Q˨�����&�Z�B��А�8��t�Oi�N��;*�d7x��e:P�-Mt�NM��{���j?��)3;/(i�?y�5�`����cG��/�N�ߔ�����������(��L��/R��{�fݡ9j�K(�E�l{�l3GZQ�MO���V���ޒ�4��m�&lWH�'�@^&��82��j�bK�j�_�:l`�}�LX�o��жFb�����1�ø�*�Q"�ܢpH���]����t�rԄ�3�M��.!y�c���|8��:�F��^�m��k�f;��hf�̶p)u��xz�BV	���ɘ,��稾q�b����COݠ�k�t8�/�o�	���p��	�ey��,!�<��lK(��n"�<�%q�G���w�0��뗷��B=a����&F�0RSN��Wo~+��L��|J\c�󒎶U�_��|�>F���G��CY�t����_�$1 �ŗ�<�Ά�zwv���lE�oә��K [��t4�����;�'n�\EJ����hҺ��8�Lcu��/�K����+�/�v�K^��D�W��X?��Ć	����Ǣ���PDl�Q�uh��r�i���Ž�,��
�U\E�3ZW�[O��*�͜r����0+L���0�����l�-�w-�LB�>Vp��y�|5h���Օ�6��e8>W��rQ�]]����ˊ�rf9򛳑�OJ,��y�$Fg�Rw.�� X�a̧�4&r�cC�uF���*M1�Q}@�ٵ�@
0���S#E�"ٻ�x�O�������+�$a5�p���,�j��6JҔ�ÚGӍ�A�V��ۛ(R'�4�k����{�RZ�m� f���R�fUl
h$T�+j�E{�kc��@)l��mH���`i��n�{�.��ع&�a|} c��M�Hˌv+�'�"��װ�pxOۍ�&9 o�O��l�W���H˽�0�`m8��*�-Kq�3���W�0]�G�����/r��1�L�+�?�tVTۈ�ӹ��}�]��<�G�Y�A[M��{�܀w�}�����8R2�^=��ͅa�_�԰7�H&��r��
̶�-�y��(YW�ɮ � ������^Um�s�ƌ���@�LB��_�A�/�tİ#�;O��lÑ�7�h�2�����g�uQ�dk?0��CB��\o���6\,Տ�z8��F@zƞo>�� SUC��P�I���E��Qp��2��p�h	�U���EC,�8�NK�;p� ��8c�	�ǂ�;�[!�N���b�����_��!���
A�h��j���1�<��l`v�j�؂�첸ON�G�@���%�.�*�P~�9X���,Ԕi�댣���_-�o6���R7#|W8�<�n��1��1��h$���3��`�6��|�x5����Y30:��'a���C����/Fp��8�1r*F��P��H"�$�q+��[�9���9�Q-���H�?�^�g�Us�&`?]M^�E?oQ��m��I�{��Y��ȣ�{�$P�4���(|�XB^n������*őu�x�?�g��,xD�]:TGS�e68p� �w}�q�sJ�w�s)-)�4��2��ֳ�]������a�h��qi'c����.b� Ӎ_X�}�aC��-⾖j+ ;���@ R�YP/��W�k�}���B��n �qdo�e��讻�Wph\fq���1��1��? B�Y�������w������H(@�ߵ�0�B`q�Ztf�s����s�;����1/��WR���Һ� �3(��e�K��[��KN�SB,<l��Q�[o��5��O�zR�����ze�SBʓ���c��\�k�7�I-'���^�Sg���Ɓ�0�@l��C�j+�Ex���Z��u=�Ob^�LQ0�v�Ј���)}�I9I�b�p�*���o�D����˨
G���Y��?���yӒCW����+��a���P�7������s�R��f��d+��̿J�=!M��Q8�G9	����x�W��N!�7/��y�
i@EG�]|��Mu^/�g�+È3�:J!m�<�I׺w�5����NO���������h>�چ��Z���.x�2��@@}Tp���/��U��h^[zI�`�S�RF&��3�(U�Y�8�X:q�3t��L���$����R�i���c��x�Gn�J�mgfmL�S(]'M�_�짏�Bt���$����+p�`�x���p>-�/H�H�����(NT���S0�z/
���s�H��	�)a�֔ذaWP��:���N��3�i�+����jj�I\MX]��%W�(F�Ӏי���M9u+C�D�S�B���3�+�J��i�����t����(��*���싴.%\^���q�N*�:�'&��q�rh25C ����1�/㤡Z�fOq�_��<��J%R����?��tǃ\��$��i�(LI�<�e6���q�"��m&������#3�p�ס(�Ω-K�Mjnw�ް���(ռܔ��(���A��U��$n�$3*���K�� � E�?���e���j��Dp�*�n��k�O^�p^ݿ~�w>�⃣�>����>o�=Z%"�إ��0����lO$�<:]X)���r.�rYM��a7�7Q\,L��x��^��u ��B�P?h��w��T����d�xn[��I��;�2 �
�;Q+�<�}�� ��n��ȁ{`�~hH��ck3l[\��d����BW� C���5}�������_ݮ�`7��yVT�.D�[9���(w��bL%�u�᭍\���o�;�Y�?�h���1E����d=��=�H�V����{��|��}�OUI�8�iNU0����N޻D�å�y�C�⏟���A�4��W�O�)p9�s[���i�О-���w��{�O��i�G�Z�
å~��dTT�I>�V�1Rl�.�_оu�ݞ
ig6ڶkZQ��Z0���Z��:4��c�7y6ʶ3����pMe?@;�Qc���R�&�S�