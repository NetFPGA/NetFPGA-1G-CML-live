XlxV64EB    187b     8e0�p����<|㓶q�P��J�Y�h
qCg��.����9ڇڶL�Ѱy�݃�z�l�Hg*?���.;[�"X��#��D�S�95*+�`"-=�xǷ��:W���~�k�
 �_NR�=Q'
zq[SUޞl�x�c�H2[[t��џ�P�Uy�Ia�T�j�9=���l�X�F"�?x+
��5�]�ϴc�2�F��>��C��p���e����,8��,
jy�����)#��[�F	���g*�TXg]�K�*�Ӆg-�P�G��]�WAH$l�����UV�Fg�^�-a��Zd��Y������(�$1Bx��DX�g�g��̽��ϴf%�������r��V+�u���./9������gn�(n��ƭ�u���h��D�R��6�"��|(f�}l���d�{�����7#�f*�p4���x
"�"̑:�!��1��w��	��bf�m��q��0�x��U���ZM?��4zH�+�B���>��YM��|���2d�e^�e�A��V��{͈ M���L�W�o58��=xEO|�x�-��z�6�%d�|/4���d?O/�n�����]w�����A��fU:3������M�7u_��sd�W�޻ֹP�~������I4�b�}�s��琁�Gd%>%i�9���G��0���;�δY8��U��V�Vf�|ӟ~aec��~2�2́L��(��.�`Mѵ�O����M:y�B�xS�'�Ocy�@}Wx���������yXH*L�����YHvu����"#��6:����ܹ_6?N����Sn���Sn �VB���0!�Z����U���Å��e���+���;/�P���?��"���$��\#�ɴZ�a��t�d�`9��>��8�J�����d�W���79z�5w�r�~��Q�`���k�<xx�|\��r�n�n{'a���*��&�;��n5+F�gm��M	�~�����V�L'�d/	�E��/o)E}RXKU6
�v��U���ݘ=���c-��$�}�X���vt��Ҧ��h���ǥ����锧�|�o�su�ZB)19��E�r)�޽��Q}���i�H"#$�O��]vL��S�$\ARH0�i�o�Ռ�8��.P��]�m��E�;�jxW����R��J��	���G�v�k�雐f��B_<aX��Ό�d�5P罬�ng]��%�Qe�rj0Z��}�0��x���	u0����Wg��Q���5eq�?�ԧ��[�Y%~�/zj6|}���Y�h��%]���Ε3�AѱS�dޓ�mU��z�J�Rv����X��#'!#�\�\h7��H1���K�L�~꜑��G��B^�Ѣ�MN(��mT��rd8ʇF�ex%ԕ���HQ��ruU%����P֫�V�<����ߊ/7����(xb�+k�۸�yzXi��L	�O���3ٸo4�v����ax�|��6�����̸*,M|�1!�mY6zgv̞���<�W��k`7�Yk�y���%�E?�}��W�Ev�D�amQws� ���:�)t����-�Ӑ�[��K�r�N��<oM��8������c�������9�L�}a�~���ȅ�#y�nr3z�G��!���8�;�]S���C$8�kJ����)��_a�i6E�|��b$��B9�GU�E=���Rr+���
�PAK(�� +��B�͙�]VE1��KV�c�7���P�
�u�uk�O�٦A�j�%i_���Yk�
�)<$~�	�\�:�T�2���R�he9���<g^U_8y�����w˝o�:o�Jl�0��G	��`A���+��i�&݅S�a�T���J˩�߮)�ކQ0m�e�vf4`�i/(z8�&�������+vK5��'��d��~�kvih���>�ݓ
�)�d-3���0yej��T�`c@��8=����^���(�C�s.>��?;vEV���%]tvɴ[�����Ar���?�!��+�\&6��:� Ni�h�Cد{J�U���E��-v�n�Ug]���@3����8��)T{�)�����o���Oo/��u�س���
�1S5=R���B�(��W7�(2�!�I@��}Ћ�Mab�UesG�C�jv����~��������f^��(쑺���kH3��1̏����^`�\�ж] �	�"%3�W�R&ŏ}�Q&)�Z0��P�t�