XlxV64EB    19ba     9c0�A�;��ʽ���v-ĹI����_���? /�ID��5"m��UN^�A��<��Y3�Ӆ����mwݏ�t��%%>�V�C��l�+9��%�Ub���@�.����e����B4�P)P��9]�!�!�����(�)O�UaCG���vPk��	=G����a�'����=f`�;N�<�$�=�,`Ij�_��7�Ĳ��s7;�:�+�F�qM6�AD�����NC1<���� !�k��LoR��	N{1�����I`W���4�2�7$^����~��O�iP��+�F�����v��Mv܂O^i��W��۩ v�_�S�`��{�&M�Ŷv�{棐&̈���y�E�8�J��f!��3X%n���88�5)�}O�):��(��7�d���V.��S$K�0rθ�~dXb�X�B]�*���79���W��`S2?��'
	���z'j��	�S˫�,x�����d�n�m'����(?������Nw�#�Ζl�P�snxs�(rU�>ǭS0�|����P��o7ڗ��u�)q�#W(�i��4yz�Q���p��L΂�B�L�A�چJu�3�9hB��(�8���9���Fq�C�1?Ì����ގG}/Q�c��)P���U���J7&�g�.5��O����IR��u�"wosҨ��H?q�� |W$Vl���#����H�D�S5A���e��`�|ab��ԕ�I����ķ`�06q�ܸX�2)G\:g��9PgI����p��o���6:W���O��J���a�;�r���vvjK²�fNW�~���h�h]�������Z�dp1\��(���y�y��!an��c~�
O  JF�2K�����.��=�[���F �Ѿ{wJ��/(���Kq�i������FT�ń쎵�g�yl�~T�he���:���coo������	!2�����!=0k��0���HKu|�[m�\L�$g�a�]���޹#�Lg���,���v9R�C}j��wb/���4*���tQ��?:۳;*n�)Ao���
��p���1���-=-�d`"Pj��T5�C	H���:��>���a{.eu�J6�H�~9��y4���$T����V�������4�����>N����&V+0��SJo���y�:m��qu)P-�|	���u�g����F�J���4�~��@��J=�?����d�,w<������^��E�e�U̴h�(I�F��р�?�Y:V��o5Y9*�*Ƈhz�rL4)��xG�Wz�'J�f��!踈���H�y��� ރeF��+Z�v��rr�[�Zɒq$M+Q���U�$Ե%3��!�`j6�5�B�xmô��5� ��~�^VzB�Q&>�KA�c�!�P��ޏ�\@�A��x� 0c(&�cu�\�K�$d��X�dryS����Ƨ
����b�v C���1E��I.Vx�H���?���|��6T[d�O5����9��.����c�Sr�U�(���4_N^^$vHYfoy6FgNZ���ȔY�Ћp����Φ��`��:�a�������n�$��ιZńP���:c�7$�
�o��(4��ƿ�<�{�½�S���Ѐ�n�Jж�-_�_F�Q�~0�끈>�;�8j���phw��3�BL?f�����2��A�)B���":����O��ax��.�k��ge��a��y�����zl���?�h]fj틄F���ʓ+T`R[A�Tw��K���ޞ�������!��:�А����x�K������4�����B1Oa�����آɩoPl��� ��VΡݡ�Bp& �w��d���lH�n�D��L6H��]�<h�02��T튮�)�B*��oY�h�yC���A����4��D�qam*&��+�6L�zI\��дu�n��5=�W�O��{4�mǔXY-Y���M��G�.*�^Jnd�e`�$���I؛��V���Je�����G�=2�r4���9i�և:p�����,��T7g#^��AI �i�vc1�	k~BL�y���zNF��Ur},ʲ���x7�Ky{f!\��r�2 :
����/���@�E7���p�QC�M�;NuQ�Kf)KC�v���m���W��:I�)��iފ��tԦ�}㑁�-�{q��^���<zK�E�Y��3�]�����N�C���?�m�\H��@Qgl������bbefk��Ur��C�}�ZV�@Q�s#Օ�
^�'�u�4~+�.��r�C�/FO�S���O��4;�[m�����r�cu-���0�*��C��;<���� �A�`ޜG�q���]M)U՜���z���<� �Q0�
5�|Z#�60w��������{����� �R���������m�S��Y3�)�gh.I4f�`濇u�;�M�w O��Ƥ���o�.�v/�Ȋ\޲����J�ʬ�F7+xA! 
���z@��)�L#z�s�ГA]��v���