XlxV64EB    fa00    2f80�bqeH�YC�%����%?$�^�h��;��OG��`��1ھ��14������I�98��lq�y�L�/� L�ui��4���P���
W�F��2�F�ɨ��r�9ni��솛4�F(Bs�Eg��5��>=��Ћt�sg�Q�� 8���~u���bFs�l{�&�"��4�ye��xF����}�T���An�sѲ|,ץ5���3�\�4/1%��%!I�����M�w�'��Sg{���{m�d��3��q��|��
�s�ru�e�<�p��c7ƾ��nXU>y�.�81y/��\fY }�d�u�V^c��&��]a�}��I�	�2G�SsM�)�d��]�ރ¹R·4kt����Ζ��G2���C�����
�G�F[B�1*�>sr�R�1�7R��U���⬦v7���Z���5\d��S!�+1
ݯ ��@��s+�+&0�-3���>��JV��6:UG�OkL 9��Cۭx9�E�Z'�Bζ+R+Os]ez Ѥ���)���v��~��m���+�ӰCG�jJ�"��[e�Vxf���]��hR�K2���.��3ܟ|P���&̳��è��<����| ���Q7�5��.��ũ�_o��qO@yΚdL�<1fE����p��#�(��� �(uw��%e�
���q��Ra=��7k���>��A� �R+N�"��LUAZ�9bVZx �̗e� 6m��[��|?1�L��9�p9��ĩ�cs蜝�BH���q��!��W�D��Fuм��0�V�g�P t�!�J_�|� ƴ<����if��F_�����	4��#.J��sb�*����}�3��Y�R�8$��bXD��k�t�i*��E��w6�}3�����K��Saݛ�I �~
q�=�Hq�P0�5�3/|��UW�
)G�|�l���f�Gh���I�wtڒ���O�\J��f�����iE��)'����IH���.���z<'������|�N�_�&(w��v�
�1�%雕0s�6�� 
r<���I��]����Ǚ�F���Ӑ��?äd��?{�p�Iv24G��@��É%ZN׊�4�5��[VAD�B�!Vu�n
�q�a���a�_B�Ҥ�BE芋�ن��Gu6�ފ�	Ji��#n���!�K�ϐ�@�WKJ���+<�G��)�
����o���-������)�Fr����o&��=�:2��B��j;�\G|�P hEW�&�X;Q�������Z���
ՁFk�t?U���D����ͤL�jڋ,Ɲ���k�n� 7xٶD��2 Mͭ�v^��b�|�:�Q�1�	�"�$�i�Ғ��_�7��Y�o���e���hi��iQ���6ԩ�ATS^�V-� ��N����n�n#,�R�&F#�xr���ʤ�X-C�R�jY@��Q�u�,�w8�%�p�w�f^&7�C"*q�G&S�)ZX�PG^mu�A�������(���<�1��
��Y�bm��65���*�"o>��'�7T&��|
+%袜��m:���O�Y��z�w֖S�]mS���ǋ�����8hl�R�D4�%+���[ȭY�e��*-oQv(A!Z|ag��j��)�� ��dcNn0��r[�-)�����pB7���ecŠ�s�ok��2��`�KR�Y(펷�NK~)hJ�� |���WϢ�+��aJ80\E���)Ŭ[:�y�ؾ�+�&�$/���?o��e��b8��h�T�Z5|�M�����
"��c�G�Mv���2q��ɭ��v��ѱw(`��V�8��.��$O���o㽏�/c�?�'�vd�;���X�^Re�F�V��'�O��>N|8��Y��z*Ƶ[ޙ����Q��Upf�5�z���O�6��,��G�X��x/W}��"��Z%S�K�=vI[<�d�֫:P�B��0�o�Jde��\�䍲l��l�	���f��A�6����LY#�
_��O?�%C�Ņ����ً�����7���4�Z ��jGi������)����#���(�ߓ��N:ZE��q^�5;
��ώ�צ���r�'���Ð׭�CX��@�%�~��+�G�6��A��	Ye� �8���	sx�ݾU�!��A+fU+�@x�,�Q�s(�eX��k�&�^kF9^�����m}��-9�r�ի�6��M<�'�C\0/V�jU��[��mo-Z�3@ᠽ�2������$�5��>y����_k�E��i�c��0�P��.�0�)�r��( �V�C����@-��A=�Kyj@���0'Za����GP&e���{��O9`Rb� {����6(H�pl��AR�Qy��3�ȣs�R�̨����nz���uP#f
O5��>�Ɣ9����3��6���MѽG��L^inG��Ci������ه�^`#J6�Mn��x xF��W������բ�����F-_���J��X ۵2�4RY�_yT�f^��}�U5s��0�To�w�� �1S�����f��sǛPq�|�B,e��m�̀)à��Qw(X������n�]VC�n�j4�����
4��~����5�j"�-2=Cp�w�(�xq����5�����k_�� 1�fgM ��Be���W������0�A[�k�6?dY�ďd�u��y����],#*ph��1yD]��9�r�r���{�H|9-��t$��Kr�M[�t� co�|�>8v�3^�xB�h�e���*�� ��#,x�ȼUm\*�Za����c�.;�S�hզwP���E�M��Otcz�&T��,�lX@\
��4=l·p�c����]��k&�3�W����F8ɉ��Ն`O�NNԾ����G�8�EA-5�=SI�����A�W��p_��>����.�8&����� {S[�Ӎ\���R�3��^�'����P�7���M�F./�w�	�`��O���K�k��M������vQ��ߊF��v�tBzl�M�Yw�u�,������Y�$��3f@�~ o���{t�����(�71kEO�vk�>��Թf�|�R��sca��r�T5�h��ZCpq�=C@Ó:����k��y2���U�k����ƶ�{��Y.��6�OT@�O�����S��%�G5�_�"�����*�}�FL����o_h�A��F�v����Z�A�8G&���І#���'��N5��a�-h��)���j��U?��¬d���9J�=8|��9@5]���{��m�*r����}+�&[(�Wȣ��Ga���(�[g}�8bDTī=�SjA<`�6��ӬG.�]���7���Up��82N���v�o��+�U����TE�g����i>����ռ�D J�02J��!���6n,�_&�Z� ��6a'��\�w��~^�����P���t�`'xL��#1��<	
96��a��i7�@C�H��9�I!�(J�C�]ׄG�h��x�"͕��C��|}�e���3[�N����g*)t�/�|�����Gho �e[-*��]��� e�?�A��I����=�P"�b~���g�O��(~-�������>�Ǜ[Ј�(�����Y[~*���%��Up%�_��w<����O=���O�*� ���4`��LY��6�}L���YO�i:7��� @���rYv�J��������ؖc�=���p�_�#���$S��_�ʘfl��8�ς�cDS�Tx�(l;�}#F��&sLS&�!*%(ڢk��I���	De�Th�MG�xW�w�5�f٬G#ĹOq%2���^�rD������G/�����k�� !F�A�8�
ʤ���2���ص�'�b!xk��<q�"���X8ƣ_%�T(-��y:������J�K��B{6PY�1�����Oٰ)V} M���g�_�Q��RF��������5�k�Qm%���\����zk#�a�0} �y��%X
��te[m����7R��j�E���!.f[r=�a~���;�0��d$���C�Y�9D>�e��Ou>�7�ևtP&��͒X��2��Z�kF�[[�W�V� ���T:�{bs��+��0g�]m;���ߢZ/4����v�t�B18)V��N�,򞹼HT���N�ꎗ�J�E*����?�I�(˕��:B�k]�1�gc a�Ja�  �ASTb��`�(L"_���Ω4������FN�q|�g&�0��o�g�
EL�H��t�F�"�~�u��Q3^<r�WC�27l��!�r����S�oV���d�a�>J��LC0tt��m
u�A�P�{]�"�z�,4�݋O�0�������Z����+�]}4�f�L���ىи�n}��&xs��q�=#S�CNQ��b[U���kG��[���k�:��Ï91����L�(�\�W�3gT�bC����%���?]8)4G'w��:u�MY�ɞ`lbT�Li�ɫK�Cl�+`���J�|}�&�$Zzꙩ�T��B�$J�xi��~*�$��<��"�aoq�y$fS������Qw~�z;�/��4^} �m��V��cZ��^�xw���_��&��=4a'����(�^#g�q�j�[�Q�����'w ���۰��21�Z���O�,����М��vslTOנ�,~�cϜ�OVd���$4���c�ڮ�5ൔG�|OH�3��L�c<M*�*,�hVC��'_�r��ґ�����gs̅�L�!L�����������7�t?���$^�c�,s�'�����m���/<c�"������v���rj���ys.Ͷd��2�I��3ezV9-�L�n�y�¥���]�����|��^�t��c:�J��6�:.nix��F�+��>�=(Y+���!����ܶ��~u��T���g�É�9��G� ��P#+<k���nǁs!�y��^��J���������`����u���,oa��\�썝�.Y�l�ᦋ�)M] ��5�t�cKc�	G��~g��:A{lV�=�NE'��$���^����"��9�!�ݎoG��H4���N�M���Gv�a����Mt�FUb��HLެ�m��S�K�FWE=$���G�2bv��ެ	W��Q�/�zo���R{#��������d�ii�T�?DB��UE*6/�6�7�z�*��!�f�˵z�{�T��[ٙt4IiZ�D}��ޞ�7��.�d5���M�1lP���֑��"h�aJhA8~1"���ً\{��f)*�n��"u�p����4�)��1���8����F����٬6����[�q��~a��P����knÚ'�� P%JҺ�p-�|��M&�s0��ܞȞ_#���I@������-�J��:�t�߸�'������y(�۫vٜ��c��a�z2������t�Ԋ6���hG/U��I�v]��I����oO$֝O��8$��iأ��������cu�vC��	tvK�RnM��b���lk	1b�C)��0��7Y>"�wP�*r����!�i%(�L�� 	��Z!��f֗#~`.�U{�A��$�!�Zǰ�x^��U������~��g��KY���~>��X\X��Q$�ۓ͠fR�k��/��Dx�����Bֳ]lWC����s�g�,֔�]��=F�k�$a�쯄,�%��|?�E�N��K�$�9�nb�HΒ١I�t"\��uإ.m��p�����3��Ѫ_��5#����=T��B�n2(��E�s�ח*qI}��D���1����_��b4�J�m�W���� K��yp�g�Vq�)�H�Ɖ`{���rp��l�"��L�0Uƿbx%�:c���S��E���T˓�9޲��Iak�����,:�)3�������|[���z�5�����G/�}!���7r�����8)L@���4W4�(:f�h���"���^�޲^!��T���';2���Z�^ZY��ڝ�¸E�#P�!F6r��� 7�)Y��k�ô3Gd��ˆ�^����q�ދ�譵���. ��0�sYf�7;bt�`�;�K~є�=Y���`�80W��"���ur���@��#��B���O �����tz%Ô(6�M�@C!t�bLn=&�����ڻ�-��k��hE@��rO�[n�A��T2pEN�L/\IЪ�������;E;�zh܈ܸx Y��%%��,��cO�e�H�J>�co�p���p\���|�m?�R+:�A��u�5�D`�{��6�G���~+�w�e �^ڥP$��td7Z~ǓA��?*{I5��/kW�����/�,w���M��6�c}4�<�DN=���8�L�l1��ǚ7�3�1��G=�����H"&N9��G�W(�8�
��l�[���*� ��q+����O�����3�H�>eV.�_$2�F��Z��m�)�X��-"E�3w��"Ai%���ft@��i��Y�5o�9[�-��'ܜSz�c6�*L�C�]U�e�"B^�����ͮy�� ��ȲͩM�&~Y�K]���6�Ӓ�:t�%�=�%���{G�g���,aN�W�/���\}����vݩ�VrLy&]ag�~�x��:V�C5�:ot��B��/2�s�i_���ܽ�]�l����i?��������5p����%h��`U��@I���+D������Vͺw�&�i�f�֊r�lނv��gZ��0f�(v@��8��v��Jvz����4�iu���:�g� L�z�Q��x#����4���5����m̙oo(�m�Q�9{B�6�~o%HrԎJ��3"@$���hD�@)u�#�&|�X(����Q;:L�a-�f�3����I'v&���5�W�p�%t����2K���m���9����ʴ6}������S'@ّ�3v�����GO�Њ�s�̦b#%�η_zV�T#ȶ���!��v��O�Z*���[�
��5�'�� �Mʊ����	�\q-]�z��� �ev��B�U�:j��B#R��%����h�{�Rf��ݼs�b&��B_:�hܟv>-֥�WS;�g�z{zvA��������܆�}�P"Ҩ���l����œ�Z���;�~Ѿ��'�7�3��+:O�"�G1�z��,��*ݏ�V��2Z5���L��jU*_������B�*5?T�-n�R�����,o��IbY��Q�8���r�$\bξ��W�� mq, r/30�8�T�@s/��;�"���	�$��tQ���u�J��ʦr�p%<�Yfq�����h���-��+`+�:���M{���3��
<�T�@ԥ=��k�<��G�{�z��ۭ
w�!���p}W��y�X�ZTHş��������AlVA$_~ǽS@��-��.{nP��7�h�pjzˬ�2��p}@WpJj�n�0"z����@�Ak��N���}Q��,I����ZI�U��b���v~�{���[�B'�Q6>n��$���vDIv�}Z5j����d��C�D@9�n��p��[�@����j��\���r;�P�+�ٙK	h55�v���.7,�I׭�.��w{Kn�F�PB��=ʼ�H?��,|h��8t)B�����=)�>�;�,��a !;���R�}��^�OXդ4%d��n�ց%�1�r_�
x�t���S��L�Sd�i�vr(We�f\-�/{	�5��"L����>���S�=�o��d��N}ʁ�ls��K����x��SƓq@�7!1���ཧr�Z����as�U��m���7@�X�?��������1���>��Π�sD�[��͍۳e�p�?"8�l����!��|�\�s�5��7�����F8����yk�tw�Z�]�z4�2���is|�ʗ��)�kNچ�hȆa!2܏�K�j�c�<��z?3��|���Z�f�̄?,3��z{���q�Ҷ��n�-��q��m�����ʪ�
��+���pc�� ']y�n���C���Rg�)�0�?N)�T��b�a=��� �Q�~�;iSq(9�}�A��/'�I���L�6�ue��G�.�K�+q�(���?~�K�5"ju�U��������T7�H����E���
됃��!���*gį�H�����1ʀ�4N𩎺w��p�ц8Hz�o|c�|)Q�{��N>&��� QM("���ǊX����:}L-����\r�&�A=��x���&��yI�ǐ�~��~���h[���1��%��A%����`�߈jS����h<�v��=�MQi�.�8��N�'�����𚟹,�&BY�#/Y)`Ν����ܝ�L�]�f_����_�: +-\�b"R���#�����5�d�en����ʅ��=��+kR�Ϡ���<8�7,�������s{�jk}���w��(E�e�J���zl>~:�zDR�ckޡgb��DJ�|W[K�T�]�/R�3��I!:褍b�x6�#Dt��Ӻ��5\o�G��1���O���	��^����b&a���f�W�����W���f��2�_Ev��qn8�OGء"]�D���
�5�d�|Q��W��� �+��DMx-/õ݇x�C�����yX0�Sބ��f�Z��7:4/6]�UMM��nz���3�x5����8~ce��Eh���m��T���Z�\�D���p@\���_s~<	�g�g�\�����5~��?2J�E�9��H�[Le�S������G%��8�����w�X<�>�W��h���}�%j�<Í=hÜQ��`n�G*��b��`~��-2�BMŶ�iw �T���\��WK�v�N&�ғ1`�༑�JY\p��r
O�ɪb#�kC:�%���-�Ά�)�����D�o�������}���uՂ�_��K���: ��TB��M�	�*0���·�ey8����߻	:��#gU¡-J!S�D��&s`j��;�J�V�T��e��
�|Od�a�֜�C�ĀX���o|���ͯft�Qp>���%�����{����@�eI]"��7���A��~�Mu�s��ޢ'���C^��a �1v���Iu�-Q�]p�5�E/��@o��щ�sR�(4ZB�-�w��P�$	���S*�o��}�X�=��q����JM��I&�;<�%h�6�3Wb�ޮ�������#/�"��Ǚ�
K�Ͼi�XZ?���N�?ia|�)��-����Ű������}Wx�ԗ'��r��1aґ�ᾯآ��ZGWGe*%�"Kgn�p���������ٹB <Bg��c��tZ��=(L��G�հL(��N� 
430����v	y>��Xq�$����FKDEe�aA���!�,��'��D��?#�`ǜ.l� ���z+�3�w���kj1��~R������4n��2:��wվ��+�8G-���IE����#2��̾䣖Me���L�}˙��@58����d?F�?vؠ����z��N��A�8�&!'?v�\�~]R�*6?$�x�6��F��8�h��\
�%����V��ᵫJ� �.��Q/�eu27����b��.;��נ�ؚ�r�V�4l0�.F�8�:�ޑ�I�-p�����U3��a��@㌅�-�"l��O��QuHFz5��ϣh%NgMH�R�[��v`�3&>��Ɉ�+x��{w��X�^��9�-3g�
�u	���b-�dK�-�����.D^�e���+�|f����]�<��7�	����P#�p��*G�-W��XD�jG�i{� a����]���d�L�mg;s��S�@�Vk�������{Fa��T�37{*v^�U�G�N:���$7�p��YHQ,5�W>���ދM?�	���l��k� �ۈ9��(�Я�bcԗb�Un�P�t.Յ��)|����HF� hf���D���b�m�/�o�Qi��c��p1�hc�hm�g5�wH�`z& 6����o1�%p�iI?�:�=܏
j��f�71�V����H���K�R���Dh��A�!��w/�z���JR~�sDG�#@f�dLk���㖎�q�/C�����2�g��J�-ϰd���_u0 |#Hr5�X���o�q���)��"6�7�LbR�E�jC�Ӷ>dm4�]��M3�3�n]�ʉP
�/ɬ���Ś�7��jm�.3$~ݪC����6�c� �Z��]�g� [�kU��J7�������ȩX�q�9�(�gKҘ����t�p�pl���g<�E�]�.��e����p�Ě��x[��A=b9o��lLV���䫋/�1t�std�aH'�m�dm(���� �#� `��I.�]}7l�E�h�~ix���ZL��-��Q�'C����:����<��aoOUB�I	Qr93�����dQ:K�3�V�p����^��u�����p���[H�����v�3�ʙ�l���;��x�9�?�4DD��3��2ѕCW�؄K�:�;�Z��7��N~�j���&�g�'� �>��psh(�%�`���l4����z�<����N���4Q� \Tz�6	����[_���3��"֥,:t@�1�������і�������%OQ�ϊ�Ɵr	��8��8�kޅN͚�}W��
/P�R�;���.O�� �ǉ.����Q� ���(c19W��}��%�<z*�B$�����U{i�D�����&[���-u������N���%*fk��&�����\����c{4��Lsh�tV�;#�|̧&bs���[�V��������V:�|m��lۉ���k������l�P=Ir�F��Lt���q��s���<�SSH�v}*���K��ef,�g3�	�S3Z���ڠ8fM'���C�Z�/�:*��ղ+?j�KB���6I�Q�3ևv�[ʶ����@=�6�l��%A�^����i�DU@b⎤'V�)0��w���CR������?�Q�<�;�:��D�{+�d'J���S��Ԩ�e�_}@LЅ�A���y�V=�̿��~L$NG���9�hjH��N^���#�*"��YvaK��׮a �Q� 3�Mo��E�`�s��^Ty�3L�r��NMpX2ZA�����~�<��2� k~֮���%��t����V.�����vl�Ċoq�i!��������"�B@��[�����|�,�J�I�Y�!ݳ�Q:`%����H�ʆ��0�CF���rp�lY��Gj'���;�BE��o�������$�-�\��r?��B�l�c��B{�^Z<�.9���VJ��� v4B$��f ��2����\@����~L��=�6�D�P�n�׵ד]Q�}1�붞�:�n��!_u84.�=����-g�hw�'=[�jT�3p�����T�bR6��ܾg�K�z��˕h��s6r���6����K��u�~	P�Bj:�/���vt4�a���d����+W'�P�s�fL�����qHlQB���N�jo ���$TYQ]�\ ��E70sv;2#�[����v+���H�?��(��p}Ey�`&�aTt7M0/	Bo`5w!�zA��=V�`�V��ڻj����d9M�����iM:�@��;��^���+J�2:���Y$��qS����ì/��z�na��p4�[�#�	�V�b�����V�$�g�ͼ��U�����o������[��`x���f�rT��Q�-��^�_�dg�԰P@���O�(ON��`��R櫗o���h�Lѡ'f�ڷ��ի2zf��]����R�Ee��/&��%l;��=����eb�T����� @��aᔻ P�r���	������RU�,s�s�jL���v!@gnAz<��U�#�uU����MJy���vĹ�+�e0T���nkƴ[׌�J��v�ߒ��|h�
.��"�=�H��m4��w����<yu�*5��ˁ@�~����Iz��s��""+1`�0�FZ�0����ݱ�Y��d���ppxTq@�ۡ�C0V7��i~)�ţ�u�ѾcI�?������cK5��������6Hϻ=d�KF0�XlxV64EB    fa00    2b00N����[k��!�H^ ��u?(�3������e�+�ұ���J-c�'i��0m�!����˿X�2>U%m�7��.>Pd��C�.�y㜊3>��Wf��$����l�S&Į%�=�.ޛbheG2?�+ ��>�;���!{p��lE0̱��l"d��t)dY���Y�:����������}p�\O���"=A�ղ��T�v:� �����~,���0�Lqn0��6d	�_H�3��&���jwn�9���GNR���1fܥ�N�BF�0u(���^O�Iet�z�U����v�=O��a��X��V�ꫳ��H"M�{�	0~�u��wD�����ǅ�پ�bQ��w���6�Sp�$n�:R�(�C&Ӓ3�.ż~�e�}HEBy�$szP�w���G#Q��'����9��
��;!"7P�O�ŋ���H�T��u��H�kѭ�G��u=�'� A��lk|-������Q޲r�H4��^�T��>B�3*�#D3�q�q��{[	?(BQtu=���I"��L��l�[��6�5���JP�7�ç	�q;�ng�&����*)��ҖY����/|��lZ�,�����9������_���{�B��=���c{U#�Đ���Ya�:��Hx��*3k7�d���ۥ��5X^�߿Nlt�ƠGf��2�t{���_��\���t�ԝn`r^t�__�����s:�·n3ͬ�G��s�̒�v��"^\<v�'c���ؒBL4ظ���n�?��T�1��Fr�B0�I.Q8O|�W�=�7�u�7A+��.a��q�"y�+�h�_�m)��z���ʾ�����5�[B���Tc㙕��Ԝ1a܉�Q�Vr�V�T�ys��A�e�Y ��ڀ�ͣ�.����>�&#���X;�F�>��N�gc�����d}���(éY1�W!����<��K����2�I��&g�E�{�%�r��ķ����Ar�E�P"�.Ƒq�^�e���@ka�c!��y��o9�Z�ؼF'�k�#�?I�EO�������#>h�3�d�[��{��u�j!;���j-�ў5:����0�O�0�*���	���|':5������'�� ���W�t5[�{��)"wz���Y�5�sʺz���zU���Z1�{��X-7��������5z���G�]�Q���LfL����Zy�_�9��S�������f�t2ИE=����- ���E��^�Ԕ�k��Gݞ�ˆl�E�et[�����);y�'�]�V��ک�:�R�&@9�b
� Y��$�+h���j��K�}�ous�����u����e��}w�&�i�(N�L��17�w-EC̪/V��`�f[?�>f	�Ey������R(�6�e�N�Ag�ȳ�4�b�a�wZS��R����j	�q;�Z�7Y'K�4�_x�y(��}�]�� 6tݮ����A9�p�Ѫ/f՜w�	xa�q��^��9lw]�z���=�J�K������rVx`q�&���ҽ�\T��g��8��.,��yF����]���c�i��c24r�DD�Gk�Du�X6@v���f�$��ݞ��/*�9[�"���M�&�U�C����\;74
v�P�	m3ڲ�ۃzM߉�Xڤ�;�#�@�P5�0�"�G#��0\��Ɯ����O���-��u�K%ɳ�us��Y��B����t,��{�eW����R�YWʶ-{�F8Q�gp6����8:�_�.@��Ѫj�Y�;�l����@��<?�D��Eݫ0��O�A��6ߍ�M	����S�����WE��'�NiW��r�Q����S;�=���m1�&
�uSahA��6��	�M9g���bKi��ߑ�T�NT1=�n,7�	�\�^8�K�	��q��èb@��	9`Z�Rћ &Iy�����:vR�y��c���.ͅ$�7��{��1����{���Cȳ型��w�$za�q���D�C�%S�<�{Oj�c��	7�?X��Tϻ�(��T�ِ�*��֎#��pk�7O�jj4�O�=��v�F�~��Ø����U�dQ�g���(�߾����L~~-�p+��f��m��`�xF���]�cz�X;0�Z=�Wa`;Q�̯�8j2{d�������<I�RӪ�Ie��W���x����r� BU`�S�f�w��_�6����q��Y\uсц�	`�W�4.��߹�<~#���dgޠ� �������E��sRݍ$ױG�I�^�R�K9�M�b��u�Wf}#�b��ȣBzW)�:?�4ww�~��C��l/����`����8W;�
}�M�2A0ß�@���R`_�?P�R���P�����[�5��Hl�����Db	n���4��k�:t%N��J��w{d�_��?`�~�a>:���2����;��+rv�Cռ�£�0(dE4�\�+�	�~d�A%�l \iY�T˚�~�q+���U�Q���d%bvu�6�d#t!oh��d\vӿ�-I��v��]���\����ȯ�s��1B�U_>���ɢ�s��2+K]z�q���*"6�ķ��y9���<�h����8`'5�6��>nD��i_U.���� �4�v�,g̊���o��Ӹ L�Oq��uzZ�@U���3��B�!i��f�ռ#�����r3��X>i�bgMC���hϺ+�[�>lV
�ډ\ �\��턵>qػKѷ9����t��!bd�;��{�Nn}��S�3P�����Tg�����&6�t;����e@R��|k{`p|��H��T�3T>�Q����Ď I.� �\/��Ϸy���9r����`��@�ǩ�X	`��~/�"o��H�À�Uu0َ�!pG�|�$��͹'�;��b��I�����t�����m����H���������~ ��i���>���ؖN�jc�w��s�<3:�Qm�)�����f8�_� ��l�9x-/M�-ZJF�6���Z��B�N&�s�9��\����  ��}�"!�]�(�����3\�/��4�Q���2�I������cY�P���Z�k	���Fcyz�lF��gD�Q�s#�d���Ĩ�sgT�P��lI�`H��\�,�*����/椧�ih<��*�$�U�&=S �C���N��:��'<=�KF������8���}��M�ШyKjy��d*���N�EH �n'<m!����p�7)�7��X�BZ�J5�m�����m�L�&�����o~C�M��|���J('%:>�|���Ĵ_<?~�x������Zq�pwz�\���I���00��9ԑ)���|>��o.��i�ܑ���mN���e.�'ܢ����¬4y UG
��|��צb��=������i:��;���_��Z��l�|�˕cD ����{�'Yꂇ��FcD��$iə	 �ks|[aSgP6>���v<Qs���!Nw�� i�ˤP��lr�iM%<4�4��ƣ1��N���]�z*F)�giu���'�8;T�zh��}\��
�_kh��X���\yF-&���ݰ�R��+��g�ٶ���ت��.cM�6�˟niq�s���">�e�5��e3��g1LAl~�s)������d}V�[�z���>5�x��Dm4��F���I�e��,ذ�i�"��fX������a3?��"��\5f�lJQ">�.#u��,"�f~��8�������
��E#��8�G�u�9�o�B���^��
���rfB��ٿ5k�uV��L�/po�,)�dβ�T���m�xrEt���#T� Ė$m�F��d���{�^�I�h��G�9�/��;��]q�g�C��d5:�a �S~Q�wX�e����K�Tb	=��)?8Pr�S:���x�~������'��O	��@3�s���;�k�:>�$�9��b`z�aL����8=y�dyX7�C�p�'���������'Ϫ�v��$��x�Ɣ�Cc��X��_.��[۠��?#ÂY���ɉ%�1?gs삝ݾJ��.2	��*_2`q�ۮ2ET��	n�o�S�Cyqw��En��"�X�
���6@�t{ oB}�R�uX�6嘾���ܗL����^�Zz��C���ᙛ_S�`��2�p3�2������,U| ��~�=5��%�3�Y���=�-$�˓�3��Oŕ���a+Ε_gz&�^^Aߏu ���D3��T�	ˏ�ލ^	��ӵc�w���4&#� �a_5��܉ƀʢ
�Em�-".�ɿ��Lڳg�j�ٽ�B䶬Ĩعc\@1z���Y��99�3��S���t�&��ҏ�cȟ�lK``�[f>�i�k���eqŝ�5�YgC5�$�����'��r')�����0nd�����P��J�c�^m;�Z�~&��֫�r��o�uc�J O��|X�ւ�4,YZ�a=���E�V0Ҁ�6m�_^e����pz�z�{���|����-1�YЄ��Ȅw��Y���u�KM㰩P^gQU-����t�KQyN?�w�6=8��U\�R���	�Hń��rw�0A�N�3�5:�5bc︅��;|h��vӒRX݋q�1+6���%�P��!��S��T[w7��\�ޭ�*DS$F'�
�IxR��1�F�_n����chK���1��P��Z5�K0�%n�SV���P��:+�[�  �O�qhCu�@�i����N�NS��p`���J����	*�;f�
}�pרJo|�q��eT���z�;�ǳ&��X��JѶ��hv�;��̏m1^=��ܐPF���;��4�4��5���H��J�n!��,��w�8��]��g�`�j���N��k�?�Ǻ���3� �!���ʾ4��֙2w`�{�I3�?���(��q����%NVCw݂GC4�_�����.�[��E�l��������W�"Ƅ��Y�_���k���P��|0�=c����k�'r!_Y�b�qa�Q	7Ԯ��
|��� ����pk�@�h�1FO�C6������d��M%���z�����A�l��x�x��<����P�C� ��.�x�aD�E�4|R9���Tp͈���ѡ��f��ә�p?@��V�ui@Y�9�� ����R�k^em�|�@�p~mm��L=g�t���{1bAm$�T�-��l�6Q�K��?���(m91Ⱦ�Åc-/�F�� ��?��$o��f��{�w���s*Tj�sA���}'��$�ͮ�X2I�_��8ka-�����Oi�9tr�n�ڒ;�ǻ{�ni�Z�ж,]D��c��5eX�d.0��������")�֛��U�����9���$�M����mEMQ8�h��(���ڒs��~�~k�xZDz�~�߉fu�uQ|߿��X�=���65��-uRF*�e� ��Pu;v��א�m �d�+���$�󍿊�����)�Y��-m��kM	x�gI�=f�%�?Eɑ7/kqz=��O�i�zW��-j� �[6��S���p�0�w��*@;�7⊍��r'7��.����*��A����$D{ARC�X��qtx;��d�r>�)W�bg�M֗��UY��oC��)/^��b
���M�1f[u��+���ȖaH�q�*�r���g�i�c�p�1`���Eʏ���{W���ŷ�I~h��24K�.� �w�}l$�T����q�B9��:�s��pI�;�Dvz L��~h�a�椚�h�v<"�}e|���52�:W��63���'�Hr��=�納|A4&g.��#�����7��5en�a/$���0PX��#��w=_����|G�a��ؓs�Ku���Ϣ�ۊ��{�O�Sv�5�/fP����j����
��]x�^�gD�S;M*.�B���cUBT��/
$&oZ( g$Ogδ���{̦�������"򾥚�ݸPl։ͦ��;r��a3�<�����!6��J4��F>x�v�!��6���_2��F�)$K�L�XlG���>�Ze¬�qΐ>�?Z�V1�����}����tE����U; ����.|=� j�p�*��B�������Mw����ꉜ�y��:+Ǉ��"����=΀������_,Ƴ�9����w�����a��A�[�5�m�OR��WEhvI҄]w%��-^D�I"t-�j�,4���C�ם���}�EJ��ia4~�V���jR�N�m�'���5�t��|ۂ�-�Lv��_�YOT�w�T�"IeN������@82��|c�F+^�F� �gY�ű����Y҃�3k�A��h��d,-��ZFPŦ�-���1Oۼ��&�9�an��C���xx`�E^����'`;��0#uҗw���?���Ӻ���H�����X��u̟<i��Jue�v�P����b��Di�\LDQK�/�`�N����������S� Ŵ��r >|�IR+Ǎ�Ϸ���G�8�^�x/dw?������f.�%�X�l�w��^�=p5����1�>F���Kf��22��HM.tkԄI�4�QL��Bv��&d́e s}uYO�?���G�prEoD�]��f~kp�R<,l0�쀲aFm�m�hIgN�t�y{A.sj��~�I�9����'����=A{C�ʦ8g�M�}ҧ�-i��yw���x'7�z�Ca�y�/n��g8��O�ZRs�$��r�5s��տ��
�Q�_(:���gp7N��aN.��֕�p��ά��$��)�z�=,�d�vZ���3��$���2�S��EO�Ndk�w���;�!��e���y�'fkܤw�"�=��6T� ,��۸o+�`94%��$�.%�> �6&�48k���8��Q�`+�T*�J��X=&��ø�~���9Nvɸ��Bsu��*�l�L�_��2�:h��K̥]�� ո��>�RӃν?�BĨ��c!����q�D,�<��BFЋo�[\�98K�(P7Rz~���(���Q1�sm�� �%U=�sJo���N����J��t��?$<�0��Q*�r��[H�n`��
4��IJ_D�D��G+���v�,osGM�P$w�Y �-�8�<3:r>�A�f�K�M�ˈ���#0^a���0:����~57,���EcN�\�1�-�e�v�� ni�w��[j�.��F�*V��EZ]�u_��o���;�sgu| ��vf��.Q��g���{�������:M��n,�5��P�7�Ͼ���*j	��>s4�#6��Ƭ��D&�,�A�Y<]���XG�KV����s<�_�a8S�n����%SZ��wܙ2��.��'9����W�?YId�cbjؗ�2kZ\6e�,�_�ځ�nh��>z�����Dm"WB���a�\S������y�'��V�<��>W|�ws��\��*���= 8}(�K���I�z4�M؏JKr�1�@�}Z�|/���a(?$*)-�#�@��O)}���t������¹�m�d��V�5@s��x�e�m�M��S�j3��~��V?V�fn�Jeᵧ5���#7����W1ߓf]�3[)@�3�4�0�&��9�;̂Q*����M�_?p}������R��%%\@f�ˊH"�|e���t�G�Uv.�L�q9���c�@̸�{��-9qd
��W��{mg��&жf&�9��M'8ֲ!.�G��c�yko@[h���|b��=�.��j��c��\���X�߻�y�1g�彠�Mk�\�z�؜��E��s�;�_�|S+Kf[�|T�tGP��Uk$���j\<g��Ȱ�+B͡�2�V�F�j�x���¿��O�z��(ܒ/����M�t��"���n��V�=�d���];������kξG���F�p���up�qX�J�E)�F|��n� �������M1r}�����+��2g������h{3>�A����q��tn^P��HN~���`���RqSo�0�E>��}s���Eɤ0��[`��~��k%(=l �rl~j

i�s�ASu\y�$�Pf��VL�>�nm`v#<q-
<�e�S���U^�8~�%��IY�-��[�J_�Ap�He�`�.Y��C�I�&3δ����#����%P+93���ٽH>1㖊��+<+J�)��m
o `ԏ޶D�K�+xӅP�UQ��[9!�*��g�ce�����2�x�T+�K���j2%#�5��2�����'.���?P��A�}��j��!�
V�ڠɓO���#�
�p��� k�S_+��5e��J\�b���5�?�,\�%j�R|��wd^$VO�P�(����fϙ�ah60�i�u&�9�i�j���8�E?����+t1�"��^�.� Ze51Qq>����e���ë�u{o/����cT�@+n��YkG���zQ�c�jU��{��e�nKg[�s3�~a�!d<�p	�hRO��#<���q ��O��7+����'��+T��1RN��{V��O���S��N*�Ͼ��<T�b	�+��)�ՒM9�C�P���㔫-�Juk_;�go�=%Y�V�~����h�0�SL���wN�9��$����u��\���~�˻�J�hx���C���7Ni���a�`�r0�m�yt���U@�/BvFh`&�����r�lS,�S}��02�Nw|�m��V�f�$��hzhm��x��I������3�"�#�iI����Q���1#+*����جu뗝K��7:�tO�sS�e%��֭�tN�U)��\4"�m��ۆˡ�ַ�$eb�EB+<mm�p��2��N��~n��D$x��ܼ�ud���(���)p;��>p��_�-5���|���܉�Dƞ`&� 26f2���q2�v?l��.���������y���Ǻ��|����j
��}�o�B,���=��ͣ�� KY���/����fI��r򣯣�&6��mn�	�"Je��1���0T���?����!�v��~&��y�"eF�RTn�_8���'	]�R�J=�r!�*����d��
N�a\��;k��$�Np-��p�{l�ѽ�@��9�1:�O����!1ci�2>��)w�čS����rD�H�� �CY��z��J@�M	Ѐ
�M�Y0]��i&>Y�˧a4i�︌n_4*�I�5��e=���Oaa����}�1js�!�D_��@���.:Ю2�`�{{ ڼ���*T�ٸP�O%�܀�5a�����WV�a����/�mF!M�*�^}��̅ $3���^���L���ⱜfۯ�^.f�h��k��s ު���AS�#�y5U6�n���+���X�e�f�;p�pH�=��F����5��pj�.���jп��?�p��!����ͺ�'|t�bJ&���ё-}J5 +
����d��#`��Ч)�%L�����/�����R3W��!6�S�jq2R��j��$@�w��9�7ϴ�p)�wJC��Ѹ6qgo�M�zR�����բ�}^d�6�FU�.P1��V�����k�����Z�Y����
o�Mc$��-`�`����lE�I�U����/��t�R���>���-;�-
�F�=�3 &̘kk�t [⬢<U��=����t%�b,F͑��/}��i��j��s�o�c*��7�iJ�;��u��N�������vQ�C���v�3/	��+����%�g���-�~(E
m*��N%#�>i�5�d�xW*8\2���XHKgP����h�O��Z�o@��U�y_'��T��6�|���«M�+��E��Y�����.�E���[V�k=J׺E�ϯx�,Џ�������a!���1���て�+BS����ŗ�e���˨�E���'�')wy�Zv6"I�8%PJ>��(��2K�STp��JJ	f:��N6��H�,g���;�38�v�\C��GƲ��0}p�B�%>u���Xa�M��YA���M|���(`�n	�)�z቏#in!|.F1��9��.��(��4�٘�Y��K��G<&��⮾ϊ���B�8�*�U�i���뵻�S�I7�����7�6hm�`"����(��m�I0�J?k�+�6�vS�\i���L�'��SS_sЮ�-������D]+�5����ĕ?FH�����׶� ;v����k���D�xƞY��N2c԰�e9ѩ�'�#QR���4�b��d�Q���';Q�E�dH��\�����'*��ʆ@��(li*n��UZ4�u镯."'�:�A��_�o��hr����'�l��:d4U U�i�����`9���J����_�dĕ]���R�9c�M[z&؛6s�m9Tz�����A�`�aإ�eLǜp8����%$�	���&��l��R�K��T��l��@�Le���6�w�=�c���h"����*������uНvp��� �r c�xڍ+�o���l���c��h6y�8@���A�$)Q����K	����Vp�
�}M����QL�U�V��P�fA�/��nhD��ݥm<�k��	���e��)P%�J!����J��H*I�_Ey�_ccۯ�ceNo��m�B�:������ɢpl=뿍��zA�2����W�,���%��#u	i�Ka�������򨝫���h�P׈�
pf�̈d����fn�8�i�d	�(O���Q�D-���l��Dm����M����*""Ire��Ƚ<DO�
��D�|~���a1F��]�Lu�^/��u��!���(0P�d^��7��������t{��	�K����K9Kc��]`XlxV64EB    fa00    25b0k5";s��"6f�7��G��^x�**�(�Gᛜ��`E̟�D�T��Z�U'�y)���e�|	g�1�n1��ֱ�F� BS��BȒ��Lmo:ܴT
{S���8Om2d�?��Q��㿆�2��D�u��"�c��	�xT�zҧ�����"<���4�"��Ds��������(�ݷC�ԓ6p��o�o�S��N�!c�g�>`�k)��=��w>�6��� Kp�ŵґy����YIj�6�}�(ok�,VɎ��<��y8d7\3���.Ѽ�*5Z��l�������Rճn2wv�L�h�j�Q*�V.۔ר��Q31�p�.N��4\�j��7j�_��I�(�[*��
��+�E���Lvvd+Zb,e �ݢ���Q�_�=v7�
�����qN�t��Vߣ�|,�-��z�����2Zp_�G9 �
���N#�R����)j��ڵk&GQ�����i�"���"�T�p�2�S�oxi�I�1'�����L�� �d� w0GE�O3k�=�Y%ә�bZ�d��\k
	�*l5�
�A�	�\|ߍ����Lk�cD�HDC��lA��}���H�#�:_���Չ�_�z�u��ĶwY
Vrʢ0���.��"����Nc��qS')���3�22�ס����f2/�Č�֜b�7?@���ǜ�\r�g�֋�gl���j`y���	6���YjX:�!�+�'Eٞ�#�n9���e�A*׸
�[���h��AA��./M!<�Ѫ�ƪ:֙O�2X��[��{�3���w&�n@�5�2`��'l4h����3�J:U\������K�V���ab���?a���H�=��w>aiZ/5���^���C�L�����|�@�I�os#$4������ȝdQ4�����T#��bf*Wd��|�{}��u��^�`�όu��\cŠ����+�~3ŵޖ��w�����k�J���\�ra=�g������v
!u�Ǌu^v�ڎ]}�Sɪq7�a<ު�D'���q�?-�W7��>{`�<���W��5]�"sa=�'���S/RǶ��_�.��ko���2��P"c������ˬ�^3v�g$���G
�F�f�L����:U+�D�b�<��f��o�^M���b�D `��T�ᵍ0�j-�L:)U�e��OدW�I�p�-bX��
�J3�v>4tul�<�}&����Nk�t�\��lG�i��;> �f��ɷ��ف}�ϚW���Iz-��8o�A��H�珕>�8m�`on�P,�J�̦N-��ds8�ꯂ����zu��2-����m��& 5��
J��zx�_/�a���p�r6$����^T?@S����A�O?,��8[F��R1oT���̯A��۳�6�m�i� ������^�SS� p��>�Z
�Z��Z��F�A���ڇaʥC�V��	��O h�l��2F��I�:��Q��g
�k�v��+�,�1��7�jW��%''��t\�HE}I�g�������r��)z
�IK4��צ#��a��	#"��'��a�9t-l�2	���*�A��"=�ci��0�!��bNr���4�r���8ޥ��g�d -������u�
v�n��(�!�9q��X�6o���B�����1a�) �	t\2����6^͝�Z���֑B�?��s�~�:�W?�oO�Z���.���c�������$����l
�N��Xk�ީ>��уi.���0f(ګ����%O���:%D��N�9�x�n�G�g�D�S[��NG���<e�G>e���W�3����q\�Z3Xԧ�y��>�a�l��W�& E¤|6�;�Q_�'� {��g:����Vm@C|�r �N��7�^)|���j�3�ΩK�a��f]|�r�i1jc�lҌ��?s�N�K	�{��� U'���o�J.���XbH���\��	章�}u��+�����{RPG	g�ԯ���2Vl��+U� ��&<��������e�ø�4�W��� �r0��%.�~n�.�a�ӜT|�����ݬF�<;�^�5z�����A5�j��`q���2�� F�uM��I��³lž���|��2��(�mc��N�s$=Z���\'��äP�q��6�X�@&��\.�}.3�wNk�=&���y_��vlKڅ��5�0�K��p��	�zF������~U O�)�d��f����'�2��p(xz��0�N8Z��Zٓ�z��w�4�X �;�å�����Nyg���
y��ZI�M���P�n?��lfx�pو������FԎ$v���yX]�P)��߅�<{���37y�4����@*_ޔ�M+���q
g0M��k��<�� �ėVD�q]��Kt>��@�WQ}�������0�E����#-"b�${hUR���>�䁚Zv=��)�5`�ڀ	\������3�U!�W_8a�rD.._|�%�X�%�g��筧g �6-2���a�u�y���.٠�t�рs1�1��* ,�R�y�Q#�g�s<y�E��]�Zᕰ�|ra��6)h=🧺â�Bc$&� �F���?=�&v��hW���||�gԮ��K��2��Lx2�C���^��;����NӘ����2��u,���*�c��ٽ���{�$7���s���d@�B�~��7�>�2��K�A(!�Ou���2o�ڬ� ���g�n�b9g�a�d��A������g�a��s� x�\z��j�Y75����f�x�H�g�dP�a沪mfQ���sX����R_�.Yޮ4�g���2�*Y5s-��e����=x�E�ت�E�����5C��f>`}��¥
bl�a)��^x[��3\��V����_����']�c~��:�/�@ۈ9",<8s����P$�����DJ�{s�p.���qL����k���*������u�>t�K6y�����ȶ�O�@x�2��������9�P��@��h��|P����c�8{>��z�5V�vk�gg�l%�ee����v��v���X�~�x�a9�:�^���{�@���Ͽa/���D��H;<�1?�Z2����b���̸�`\,E^�R*P����t��TgLg�r���#σ�2�]�lg{xB�|�	�_����q��a�Vv3�"~'�W5�����6hmν�=� �Ԍ#7'�?�/�E�e(����9~j�7��l��yx�b#���_q�!�WO�p@��+QRB����\� �H|��m������x&�θ�R�����$  ���Ч"�n�~M����h�!yt���8�H�<�",�W����ά3@��ř����{%Ⱦ��C���RԕO�|�����CU��dK�����P)Q>�ag�+��D�Ė-�8��m�`W���,�3�D�rC?[y��r��'mV��>��J��R�ʎK��q��p�@?oͬ1�����6�|�b�����.utR_�s�Bu� �J�:̂x҉߶|�zI�Mf5�H�/2`i�`�w�̅��MW�� c�h&.N6S�+�T����H�1i�C�:6\w�|�soCm�@�-�����x�]�OV��0,�i�$x$2��M�	�8��z �fи������PR6J����d�f�F��V�K�E?���[I&�E�R1/CX�8��t�`�TD���^C�f�H�ܟ�����o▶Q���,r�n������":���z{[a/V4���R����h��h�� �1�?�7N��K�e�`$���A�\=p=��tU'���H � 8��:�^�w%�z��M�1O}�y�=���{�F����8��J����!F$=R�H�Vs��j����`nB��U�qp8���|�"�i"X��c��"�s3ƶ��z\\x+��-�d�ԶW�F�tf�8�0�U�z�����2�
�`�u�z��g~ZN�Q�"�y6"�LZ��I?�~���9��&,�ee=����p�2��X��a�S��\JCj<#YJ�oi"J�q��uXȿ��N�2��e΄�S<�H����H/�c������hs���8g�LY~��}@ib�|=�1��0��[ 8L,��NO�O��qRֳϢ"����ō���*[_�PY��)�A���l��r�
5�+�A!/����>ȡ;2�[}�;�b�}�P�1w�-���*�G��/F"�A'�^������<���9G���;u���'3�\���E)g,�t���U9���OC0
�2���c�	%��mi��w�ӻ<�DSA47�����9\)���(p��d��W�e܉�;PN�����g<��6���kG�P���8?�r�i�Mp��~t,�ö���l�&������n��&�� #qh���%�2U,�`Q��lg����iFF&�sZ��B���wI�mH��͍h��	o�j�}"զ��=���s�8m��_��x_1O*�v�FyH7r����{�H�^�7��jH]�T!��4��c����/ƇH��gY��D�8¯?�	�x#�_�D�۟�7���� �%6z�e�$w{+�֔7��.N�ʷEI��6��} �T���3c[��*�T@��Z�Qp����E��st*n�^�M�;� �5)vi�������7�]|�'1Unݨ�X�p�I�,@ti�f>;|�.�X@d�������ǌ��A��[����9ʆ�qCS3Liο�w:���Xg��Y��5,������>	|7 S��f�*�+kZ'@ #S_g�s��d_&w�$���]�9�78���&v�%l�}&��a��j�{^J��n휟
�uwSge&��%d/.5ˮv�-Tm���TU6��]\hB�r��O��}W*�}F�����WgG[D�\[��n���c��KO�m��T� �I�)n�F9������}�����,���\QU�Gfl��)A���h�I8T<����s�ٲ�M�� mQ�?���-���ckg�:�:���T�hL����o���I	N�h�T��c��~7v�D�L��᪉M�xR�S�V�3���.@OMX��W�X�mܮ���f�� ��pE�uФ���?
�2Ȩ5�%R}#��kqbZ���F/��������l��e���,w����}�3��1U�����:��x�xכ��ݠaV���z�̴���F�B���U0s4M�vu�T�Ҳ��*���m~��}L����,w�Ģ1ԗ��K�����H}�/D0_9�ˤs�P��������t�%��.�M6*QĬ�1~���B���'��PrU!ʝqaw�te�YԡC�I<ҒmF�@PO�@֗��
|f~�UO[bAV�?`$�<�� �*�PيӭOz���?or�$��B;���d<��"h7+[V�M�����z\�Ȝ��/�? ��4�,�I��B&��
�I�Sne���`î�1w�dT�͸��i��ֿ)���F���nwѽN���X&����>դA�*������ќ�}J��ip�u&�ߠM�t�|��)���N ���Cˊ�ȵ6�eU��r�ц������A�4Y֡�k�,����3v�+{�m�;����GWN��7i��@#�exj�	�ō9 VCkǬ^���H���"�S� �x\���(x,��/�oNZ��=�,�{��4�^�{G0�2dR�:>�z��c	QB�/�����.kB��M��t�Q�$*�� V�[�A%��/"+�Mそ�H�[���5*�+�:���i��K�����M�A�S�x��2S<�)��M��Db�ZI�m�kH�Q5��Q��Uo�޻�������Z Z&g�%�3�ml��H�ϖl`:?���|�c�Z�ʃ�DŢ`�HJ]�0�Q�$��3l�(L�ف�	+U� �zO��{�׺�\Yb�/�Z˺�R�#PHF=s��'p k0��Wi�^�N�*��q-�� '��S�@�Z����i酲v�t�jo >*�$+�с�h�[���x�Ч9l�UC��������e&P�55����{�5[�徲q�<� �7��Ԉ���"a� �M�Bv�
e�D�U�-�ɭ����)��v��}ǣak�Gx(�obA+�-���o�(\	�� �dI�~�����]�zOXs�q�� �6�u�s���	)}�4$���!_�WDكJ�A�1�×g��a�[��ܽq4Of�X�����͝��=��ؙ����a�ȅ]L+�%dVe���F���a�^�R#~�N���d���1򉤡���+�@O��"e�� ��G��T��E�km]���,D�c�l��P�g$�PP_�~ߡq��V�W�R�)�*\xUH),���a�N��Z/�a������fs�����䄼/������݁@���s("�li�RFh��Y�H��+�f���0���<���@�t���>J��H۪`$t�uwǾ�ɷ�H�k)H�^��i�@'��aw�/y=�$�.Q�t)����G����bs��H�s�2r�`� ��g�ɶ?��jP_��yX�WLV���B|�HJ!��w
,�g��X6�`���.�fD�VS�	��`�J�^v#�)q5�����V���� +�w�_�g��~�f�e��=���t@$�@;���@?���+�tX�">�����/]G+e���@?LL�:�϶m7��i�ᓍH\�B�C����#ӵ�I�`�ܷ.�O��C~��{}��L��`|���!=fr�t刌��u��e�4P
Y��[�Z�WR�kGwI��E��|��j�f�<�o�?&<�e�Uu.̐�㡅�"��Y�C�c'cy"��9F��Z�/���FF��Ntaz+�oܰ�d!�vKU�f�@�H���:��jʮC:�i�.�u-ጤOM��{��.W�͡M�/�V�R#��`�ZPUr�ف�Cx�qEWև�o��T1y��,T���������/�&��=��K`E']q4HMg��)q.��W���0�����y1��j�{����Mvit~y��˖d�"���y
�ss1vi<������`gx_[仈���+2߬ ��Q/�����lp�hj���1lA�"oV��jS����Z���<���ϡ��t��y|x?r�>[���!$�*��,i�"ZxTz<�Y[�e��Jt�u��Aa��<%#�����]HQ����m&��t��H�51�GJ:��7X�l3�#�;@k�>��vJ�
{�����H=�lU����h@�R��B��PU{QdI�
}�����@67Jɽ�SF�s�xp��zغL��Y/�r�������H�7��O�{���d_-|b�ӹɀ�:>~(O�s,B��<�v{H�S}�|�_M�P�i��?�ߟ[�ͅ���	0;l��?�����*U �g�r}�z��qn���w��2����D6���6�oE����b�N�̭��+�#�v�?t�]j@;��ƢZ5S;c�ٍة#�2� ��_zS��CCx�Sڵ����𣯿�O�ff�ѯ��å��U�8@�O����!	��\5��b*��%�)�n��3�@;�/�	��� v�a���Cv�6�k��� ��@^��ne�����>����! E5k��<�l���^*x�L9G�jH�����`Q�Q�[�?j���uRKh��Id�>�:�2����[��.�f��on���ɚ��|1|u�ݫg-���e����V@"1H��f>�A�
FPEAh?�B�.1���Y%/�X� a6��qʴc��<��W~��x��獶gs+��#����+���7o<W��}���M�DZ�=99kinO�Q%oS���n�r�
��uQ��]G���aYY�E���w�JT�]:%�q��L"S�w�0+�fq۟��*C� G��p�b�I�)�ֶ��l���
(�����j/�rk��5�J�ۼ(>��
C�;\hd�9s$9?9o��.aJ�������Ϳ �<���X��\���E���Xh�Fe�.�'%�;�I�����7�BOO�2%��5����ƴ�ɉx)�:/9 �%�F#�:��~������r���!cb�iA�*S������ rnZ^!F|~�KK
���]��v~���с��^d*�CUZ���e��y�x�L/zr�����k�+�	~xZ��z֋���"��ý����7�h&3,��y��0���h�u�ɷ;���e�ϸ�$8���_vz�H�Z�]��zbnѮ���!���Нw+�L��4�GF���D��{Eii���"�`�_u���Yg�]EsM(�LFCF�EҕXu4��tM&��4U����nFm~���
;���);;U����ϳ�����CW���җ��
6���F:���d�=l�Dm�(^_DQ��/��m��G1!Y�7@"^gM�@�m�'֕ϻ�"%�H��b�O
)e���Hr�9��`���9.`��d��hC�>鉼�9v1�VtR��2��έ4���}fw�Y^��t�|y���v�ދ�A�c+=YOT�<ƸDG|j��=6'���#�2��I���E�{y�w���E.D���c"�9j����NUD�sT ���Iv�A�*��UO&�-S����#̢���H�X1D�(y^���.ElU�TRQ�"�<�w78���F�En���=��H�s{9��Q��g�_��it߇rm��n��Ζk㓏�<3u6�.�s�^�	#X�*;FQ��Nt��D�V?���^�|�޴Ӛ���.�'ʞUG48)~�v,����'h���0wE
6�hM!@n�:��~��ŵ��Ҝ�CC���ٝ��9��V=���OKw�c%[�E��i�a�v�@�����N�}����	�t��IG47�L2b	��E�>,ʐ�{@���7���'��f/�,�
>���$RYI�xhj�j7yH�X�ݼ�0����z[/nZ�1�4f�?4��AMҊIfA���\��K��&�Y�8�-7\3z^��6��ٷ�.�"BMe��b.��p�=,�:��{�d��-X"��N�mc�^�9�b��n�.�vW�W%�Aɡ��+_��O�
���ܦ�a���=qDC�#�јE�ct�Y
�C���,�{&U�g��b��a�Yz�2�vB���מ3l$�˙�R���g9_i'X;�jE��I9�!@r6PpgK�������$������f+?vJ`�$�P<h�t5O���LSgx��U=�)�m�EJ�cW��d�C�ϒ-`|&n=�5�fN+EL��3�έ���2�Y��q���E��+�f��E.��FY��p�Қ ���4���q��;��NJ�b��ݿ�`�-��Xy
�|�
��k�γ);[�6��!jħ��.���pvi0�!}=����/J�)������ür}HN�V!�*R� �ѤPʧ܍z��^��91C��]EsdZxS��K;�/*v Hn�t}R%�6�.B˷O�����-c1��r�x�(��*� �o~L}2�Ӻ�����3�����zXlxV64EB    e24f    20d0�X���F`�	�%a)/��;	<%3�6g��������D$��J�b��iv��Vn�z0x%�_"��%�e�Ȇ�hV���n��Yr�i��!��������H��GY_[���|��b�N���xO�yO�H�EH�.'�W�z�C���d8'���AU���IO��,���w�V~i����Q����G蘖C�[���I�x�j��6N��+�6"�n.���,�)#�C9j�E�wZ�m
���L�P۩�h�������0���؆P�+�&7����&S�Z������Ժ �w&�z���V�1�-I�8^��/�F�j��B���:<wJ
�i>���*�������NC턼C�)8/��y\>���
�,�k&"�BԒ�5���W��2V]�0$P�{�9��[��x��,��Y����z�Z�~���P.(�{�W��bid�*b��x�/���ܻ�%� "�*��NZ�Z`�9{*�-���F��~UVS�����2��{>�-��Ψ^x�x����x
���~Ŕ�ϕ��êB���^\)5���N{��YU�,������0��χlgD]|:���;���!�|������%˸�_!-E����9.���1R��N������!y;h���l��W�[�'q:gѲ5ugNW�b!r8���v��0����ZC�D�ٍ�w����	�_�aoJ�'%׹e�?aӻ�O$5�bѺ�ؒ����ҽ�dfV���n#���M��f��W��)��Q�&.��^\�֖~^�,D�ys94����H�WX��9����<�����Ҿ�6j�C=��-�I��%iCh�D��|��˫t�&��}Y�`��?O{�G��ae�{��xg��3�� ���50���Z�-'�ޛI.��'�V01�T��N�:Ɇ(�g�.�uQz�l�/iX���t�E#Ny��X��R?�Ա��*���2����r�:�p7zL!��s,�Y��Z�5UqN��֎{���gNsAUn�o�ZГ�	K@U���/R1WJ�FH���gJ���e�r�n���?��2����ͳ�WC>:A�����	�SC���n�5�;�Ŀ�5x6���k ��kt�恮��#�GuvJX�٣'�@������6g��+#��r.+y�rNgG��#<ѠҚ���,�G����������a���;���^�=��$��B�ֵl�z�K�[�Jz��XP�g渗I�m���jz�Pl��@Qc��S�:Ʃ��)׆\}��=_U6.�9��=��))�J�\���9Z���sx��u�˛.u@�a��(���ׄvV-�T5�<c/�v� ���k��8e:�Q׋&!i+�io�<*_Ů��^(���\ �Ƙ� q{�t���"�֌彩�iL�J^`L��l��[P���ף}qN��Գ_@	L�c�s�@�������K}���h-RT}&�.��j�QD�܎�H��,0��dIG�;�� �!N7ɷ1�q�Vc�=385��dy���tt��Gݯ�Y^r�{'Y�'�����m������T�^�tJ�rvКL;����G� �W���V��辻յ�*�����)v��K2�x��>,�%�T�CI6�͚O�3�R��3[���@�p�s�4�}���[w߲<l��q`��2rQ����2�|7�֑;*tW��_�Su�)?V�B�
��e���,;ɲh���&+Z�����|�Q�h����(�!d|�{M�X�<����=��iWH9m�ا���oj:D�<���fbmj~�2�!p�L��*+�; ��a�Q��=��!��R҈޲�u���=��q~s���J��9]�\Ux؃
�m���Ų�Ƣ�ՙ ��͋�n��	�:r^s�Z��Gn0N�,��>Dy_���<'w��k����(F�j�SxUt�Y��V1X�Q<���}d�+���\�.���1��@e��?^�G���8�-�� �@U�*i�i{��X"��=טO�֤a�v��.t�=�>����&rGmlZbL	X�!�P��䶆�:H<qe���������S��&HE!��^����=�S]ڦ��"�!Y�O�R�2�h�
�6|�h�ow�V��h{e�#��k�aQT�?9����W��&93*�=��� �b|�L�<���k��o|S�B��m,J����L�vr�}�c�1E�Wfõ'�Lg�-Bm������M2 ��t&��HdΡ|�;�I�]l����������렌{�2�i���g;������)-<ݎ������D��H�^S:)@C���)V���gԾ��߰��Rپ�^])��L���B�s��Vh$�����m�k<zݲ|v\p5���藓v��}=�-3B�|U�����<����?+]f���kk�Vhp�;������Z=F��Ֆ���$L�e�%Z���e)�,����o�s�g�3�`�,��#�0-���~Ś(O���mt�`��53��	4+ʥ��S�.r�%�5�88��v�$�sU����Z��hb�E��,S��/�hc�o���� ��W��i��DO8;��K��-�a��Z�z�4��߻�hՇP�E�Zv(�P"H��4�C��aq$]�����k��C۲F� @}��T�}-�}(��jF��Ɗ�`]��������eҬ���A+��7�L�qc(�\���6>f�G����9�ې� Z.F��ϓ]M��-뗯��֪i*��=�]�g0�z \c@�Y�H�k���f �!����g��6�y%��q�%����=׋#���(��>:k�Z������>2�(g`5�2�*���ap���
 v�Tt��g���hQ���sG*���*E���E���W�Z�s�K��nL�-6a������NO�~걛hI��?��"ר���[����Lt2��A��8�ɼ�����sW6|���In^�z�Y�l�4�}�%��mC$!je���bL��Ó���a h/r;È͟�+plYJo��[^��)�
=IN#J����z�"YyY_����/-�g�l�k���(c>�>c/�C65� ��p/��<�����u?�|G�/��o5V��� #l+7HO����Zw	AY��mEَY���j�{H�v��pK�w���.�>�+R���觮 ���<�����;#jjU)V{��t�$�U���3v]���{������qÈ�b`&0�7P@k+�7����/��㞌��w~�h�rc��͢��9�`;j�|ҝ�|����&H@XQ��z0w�GTc��*w�+�I��¿��ehu�V�N� q�[���k�K�#�Y�W3� UOK�F��H��hR�n���NM2�;���R����R�Co�9�A�a���pr�;��[a	e2-qKũ���z"Ϙ��	��	~��2� ��%/v�U�C�@�{8R�އ��i�X��C���	IG&N�+��fb��Ky�������C�t�P4|��1Yd�i��\�i�x�ے=�|�}�:U�j*�}�!����<��p�|EI�1�I�g�M�tbD}[�|���X��;��d�g��A�ڮx/G?����CDZ�,f�J[Ax2C�/�ŤY�O�ޢ{YG��M@FN���~����:�7}��&8�c;�f҉����aye������Z/Ma�I��<bU��W�ӂ�N�Y��M?!���A�3�u�q,�)7� ���w��/c��b��j>�WZj"�#��0�M'�G���:c��K+x��KFI�&�����1���x�9	��S�c�IK��y���	�}�n��>��ߥ���:`'��!��f|^���>l14�i�m�hPw���#Q�p�I`EPR��<���t-�u ��z4��&I���E��j�t긥�f|�Qkt	�T�$��e���2��NR܀鴖���s
�A+�	��/�:�o���@�����@ۍ�b��]գ�N���<�)K�3FZ������(����q��>���4~B+�"��P���hʓ ���k��C(X��IQaEv	'qvFgd �;�%�7��7��E�ԯ@ޔ���M�|����V��X���>��-���V�*�VPF_J� }`�Y��)�X�d�1�G:V���MP7NB�.�za��%��T�1-FviȬ�_��W����Jbp��yG�Y	w����|m��&M����Q�Z�=/-5)�!��xΩ�(���A"'��v>�_�i��[)�f�0C�Ma?�xgv� B9����f[�X���(�PY�f<�t���Զ&X+�3����sL��%% Q餙"o#�!�^�� �OV�
]�7l+�hƟ�P<T��"���B6���Q~ޮ��Zv���z�`�'aN�,�MZK�{�%����7��|c���	t���]��s|*�:,����?�vl�a( 8���m�+�;Ft.����;gkQ.���'�������AC�|(�ajo��O�R���ux��۔�����>��l��I����yI�9�8��eQ���)�����?0�`�0z)��I쓞a�7"�Z\����r���H��Zx̚�������S�Q(dAWg��kX0���pH��g�#Z
=�� �r�ʟ�kæ|�o����ck&�X=p{0�=P⊟��@[�v�B6j_�"ȸ�31����R�Kk��ufy�0)�]�%�|RF�1:�e�~���G�e����t^s���h�ND$��x�ʠ�OskjIh�^4��$�\ v�f�'��8�y�g�[��,ska9�7h<�`d;K��*;���@?��^��f_����]�`,~��^ڗ�7�'H�=�JfE�5u�L�ߨ�1E��N5��m#YD�ݩJ�����\
��\7�{�s-�w����]t���4�d��������m ԕG�(�%}ݼ�!u��C�f"�.�;�>�E����/>J����?7��A�Yp��=U{�G���W�&@�q��#gc<�4ZS�#�0Zw�A�R�� L��P�_�$?�+ ՒA�cR!����1���?�fh1x�4p�~.W��I�a�ÞbG�#���eH/Yjo�AI���xJָT �cow���ޣg�B��Dh��	B4�ԋp�fP����=�-��K<jl[�S�*s�˾����$H�D�m6��(q�޿"_&��l��,�:!�-NV��B��q�-�`�t��`�7d�8����|�
6�K}:�.- �Zv4�)y�!|�����Øɯ6�u�U��Nr���FC����x1�&&��Jǐ��2>RN�(�%�}҆��=?�ej�8��,��7���	/�9���̬U%��v��1�w�E
����%�K����3����p�2�oM�:��m#^6��o0�M���J$ʂ�?Ҟi���ҏr�ݝʖM�DkD#�t�jqKK�8��t�LN�����M5�wN���d��X����b�!'K��0dɈ�q\������N�Ʉ����*]��;:��Bф�_�X�n���sS�ع�h�s�N�e^��?��ض���x��vR�,Ws&�/�0b���J�� ��f����n:ʹ�^��t�)���HjA${{(K{���"�Á���M�'e��<�n��X|���εQ����NB��"�� S�b�9�{��c}�׌��B�+���#�wTlSώ��r�a�#�154��T��m+
�#}�:Pפ�����.����������n���=&�Od�6�RF��3�o�ץ4�\��<�'=�.!����1�Ԋ�R�%��,s�_�:"P�5vL�7u�������.�`������IO�,8�Ӓ��~pl�6nȒ��O��ss
����G7j�-r¢8ǚ`'/^I����w*TSP����]46�����q���+��/5��b����h��e �À�k�ȶ�/a�Fu�ij��d�F��S��Uu]��~�k�qyE��{	ڃSOu�=�8�y!�%����T-��ۊ��[����	nAl8�v�3{2����L��H?�ߧiD��w�J��^�X���k�8&��e�z[7_c�^a�S���{�f\}�)����}�>��hp4	IthI�
��1�C��d��� |�ٹאj��M�>��C6��s��xR�,�a=3T��g�s���3<�T��bo�㩧,��(4���L��/Y0�t�pC�S8�#�B0��/��!���ێ�E�3������r�RlU���o;�_���l��f�qzMkH�P7�As(u��Nv4]���<�o�N��:��v99?l��.d�/5�o9a�w�P,�5�ғ+��r�	o/`c,s��-�h^� �Q|��q|!� �m�1����<���<R�!�^���C�t+���/�`�HT�t]g�=A�L���$a�8���"C�`ic)asR�j,��"�����b7#�7�¾�qi��b5�kj��G_�N2�5�G(E�6]@��������߃s%m��TO��&TM�G4�Z`D7����7��쾷��% �PR�+|�B{]E?@L�/���P��6�����URG�	$�r�6檂T'�թq�g� �4����2��8�w�ŐCmy1��90���]h��WC�WML��$�v�'�ǫ���� � ����
?3~�+�G�"e�f1�\�;��|]{ۄ�>�#_]&�6u��l�?=��<���cKe�5�8�(�j�ίA;���f�wN�҄�6�E;�?q��u�VX�9n��F���-�=����mKS_oȦ,<���K�yᡴgFGM�F��_�ˁ*�&��u�w��^U-)-~�����ө4�Ad��r�x��_��b)k@�O^ܕ�
�:�X�6���cm�~qk$����o�d��=JӵZ���=���ɿ6�s�O,-��7�����a�A.w�X�]�V �;����}׵U�Nu�HD�#�����J������ �3��0¶�U�*h�mٓ_K�8��2�LW2�0E��������^�l�U+AZ��ɴmUX��/�͎�ix�T��&Fsa�� � ڡ�9�c���Rne�����V���8�6\7��&y��/
�Xˋ�L�~M�1�?�,!���+����za���Y
40a	�\$,���l+St��]�a�T���Ԥ?S䙔���T��w#�K����q�%��F�*����IzW�Ɉfn������-KW�R�ah~xIj��bH�|��
����~	�7- _���y�=�I��|E`S�NSt�q�����j�7tB���V���Y~Q&�"m+Q@��n�f�;P�M������H��-�Ç�\E���n+���|]�5��U�BJ����au��ac	+�k÷��6����>�q�?"K8<�(H�,��>p\���>���epZ������Z�P��w��7.r4SR�E�(R�s������/��D����8�ܓu>�>F3ɕ��O��V{іU� �Gp8��a��轻܎���h��蛀{s��zy��ܶf��.$]�:"m��l��Z�í�?��lA-y����h�7t+������=��"ÆM�jW��3�����}q�"�������~��9�3���4�7���jQQ�s�`p��5y_@�*��xf
��/�h�
h`�Gy`�MV�M����:R-�sy1 th����#8�P����!"{�"adwaR���w�T(_Z�����������H�T��,���u�V��8�H�Q�s����Yi��%ڱ�MC�JdZJ k4�����Y>?M�Ԙ��q�	��)��,�g�q�k�z����h�M�3A�Y�J0{����`CW�ˑ|�鰠U����>O�l#� aT!�Z-�Pu6��N���a
�E^\�9Nv�r��	>"h7�k���)��^��� 2Sw����."ne�*��4X��Ӽ���z�߶����yo�+*׎kk�!:Ɲ�K ��'��~�#B�4|��/���Fg��瞜�=y��#����=�8�s�I��fN�����	P�l]Q���Eq5�.�g\d	H�:����Ψ`�1�ғ���(>>����&N��:ޔ:�X�%�j�n��pC��[p��x�s�!�AK����{2�Ϩ $v:�1,8*tq!�gL��y����T�f�̴��ݤ$�Y�z�Y.(D1
}О�<A!���/fK�0>!�<��gh��"j�h��w}]* ��b�9���#���. �\� �