XlxV64EB    53e7    1140%�g:���F��0�QVw%��ֺAj�Ah���5m�u�-E�N��_�B! �'�o��h���gOo=]0�1<+��	�*�#e*��6=E�;����ݔ�Xp���}F�;l*�\�h/�6I2�K�~��G��hh�8)'˥ �)oe�e����W���?� aF0\������mR��ζ!4�Mx�L�\�e��甛��Q���F*��1W���]g�L����.��sW���є�uh�=��[M��!���c�=��U+D���[�]G��Z�F-'!xYf�KŻ�o@Pƴ�9tH�04s\�|`�?�* �^Ӗ6�oy�7ZM��{�?1��S���O�F�֮�:U?i#�xR��Z��Y�+�L����;�����/UE�e�y��yh飲���Q�C��a���q�>����Ș�[|B^s�9-Z������a�{9q�A�H�ض���=y���`C���iJ.4�;-��p�r.�^�:�&��??՗�=��Q���Hd��Tý�f��:{J�H����j�"~J7��2W���G�)X˛6��m�xd�J�``ϒ���Z}4�Y��>�Cb���'�ۼ姘�����E�L·�!w�(��ӽ.����5����<m48�bH�<���K坷zLeޗ���|M�k7�z8���P�^*V;���%�.�75�#m!$�*)PB��ꛖ �͙)�����m|L&}\�p��'�T�%���|p��
G�'3�a�m�7Dj2�I��Yc׶���;}W4���������q.o?�7�VS>s�^�&cRza}B�9�^c?1��L*�>������nt�C�{����o�}�<v��,�XҵO�`{�|��ۈ�-k���(���3"�x_��#�}��ƚJ���Н+14��*q������vp9��i�u�V}RrbKCY�q�G?���~>la_piU<9 ���� ���9�T�!��Ò_�P=� 7�҅�C��g�X���|��d���	EG�0���o�J2m�
�O�۾ԃ��e�:�bt�;���	j�~<���j�{�1M�v84�./�}����k��X��(R�1�؇��0G$E7���HH���A�Pj���S�"��v��5q�T0�7E��r��XA����Ǿ��K�6�F���ծ�p��<ᦣ��fm��ۮ��W8'���RHok��&C��{@�޷����x�J�$���ض���Z�iRҗ�˿�bZI�s5������㣂������K��E{�y{��?��w�^&T3�m��,��Lk�C_Bo�sB�E�����Й�'B��kOD~i�SU���D����S�������.��I��B�<Mb#]�<k��9O��7�&��Efa�.#AF��"%��ӪR9�Z���p�t��@�>�j<Ot��wrR^WA��*k,|���-��d0/mp�Q7v�ocS3*����R,��	
)M�}C��R�i��r�&�ak��t�%�/JT9����?Z ڪ1;z�t]�3����U�Eɫ�k�Dǻ����6�z��^:�dW��J�o��b�S���Bġ�/�&��3��o�#@/!ra"��V[t�����i �.��"��%�"�-�:����!j-��ikC�N�F`r�����8��Wq�����u��ӌ�[��d�4	�3�+��2�n�T&&�ҔF@���JD����h��16bH��cs����55��/}} �ТV��o��&&4�1���`�U-�P)�lI<���m��*6��L�<����39E��E����C��BgM�|d܈����ˣ��$XE�;�:���+^>ս�����<���x��yx�v�mw��(��y�ש{��m�1<��3td��ނN *��ͭ��q�>d����U���Q㿲-�h��5�d����R\�j��f�ʪ��̴�ɒ[�IW�&���h�U[D�UZ���vox����`�8�E}��� e�N�>4ߠ<���+�
R�j�tx4�NsF�C�6�O��.�A
&O��2^�t-v�I���[�r5"<,��ѩ?��>�Ru^(����̑\C��-a)�I���~=A�
�����np�k�ɑ0uc�2n������/�sٗs|~"@��*��w�	CH#�YkE\*� y��(C�H�'��q�=r����F��v�宙A�xB��3DF��r���NB������ &{��f�#�i�)�@� �p�⾯Rq�/
�Y=��n\V�k;���<�]Nh�/9����b���d�>\�'&^m�����(y޼��M��V����a�+��BT�_�'�	�P9�%�;�hv�pO��W����</̜A�ׯ"3t�����+sb�l`M(�2C���92+�:���I����k{��J6�K���8��1]��BJ�Li�EU�b�X!T)�pd~���WE9�x!�p� [
�6��̌��z���N�e���1�!� !tk�����@�t~��p���m��6[��ѷ����V�{ǆ����#�]%Q��䶝=����|���9�w�]h�?��j��t�+#��h�BlL��o�$o���b�~by9���j��An|v�|��r#8��w���	��`4}1�3_����RJ��iO����|/�Άnp!}D$L<Ё5�ߟ��`0���]~��G@�]V���rƏ�R���CX1��h��(��t�1��tg����7ꌝ<	����i@պȫ�	梐�p&���@(4�9(@~+j�v�fR�fK��!1ʺÁ�A�IPyF���!�gZM6;�}	���o�d�YʛsQjt.«t�+��}md��	1V�>�7fY�����35�/��ZC���f�;�gF�P .Ca���*}�#c�W^���8��pu��+a* �	�I��5畧9Y�8(��������|Ұ��\p�?�|@^��3�6=_�rk�SUh��.S]�@*l������i���J�{gS�2S��/��n��$P�O�YRb�a�v����b�K�g	O.�J`_�;��m�K�����1G�BI�3N���*��e����{�~½�gT�-fgi	��f�f�ڪH'\u}�,�(�b����-��#��9�����eզ�ƚ�w����C�����w��C�X���:߂�zmKj(=v>�2�Y����0�z0돗( �?�EX���kkI�R0���NW�β~�o���_ �0!4]��ʬ��e1�������<�h�_|��)����k�2���S��e�U2��9�H����2D���k��#�?s��ǯ��nPԬ A2��������;�G��ڰĺh����Y0%�7��/���iGt�8��Upʀ���ђ@ߤg�߻(���bJ\����Q{�e
�WlLk��~Eai �b:���ٌ��(16U9G.NtF'/��郀�;��R���en�m�_�1@ޥ�W23���,��t����
�Nf�JʈYMR���P��s��矤s�BI�d޷p~������\-���u5�VԜ�p
S�&)�����\
 �ٻZ����9Ҹ�oFZcYd�����HfB_��o�J"QQ���oN?�ﱌ:����k��ļÎ����͆�]j�[GZ3␇�zK!�1��w�
�V��b�"-�đ-��0;h�P��mcn��L��os����Y�+n�n4����qwR+Y���y>,����ؗF��T��Ly��Zx�w
��"j���8��]���~��3߭0�m�az��N���~�i����MI`��C��+y��7U�YNѲdG�W���b�+�[�`�6���������;4�,i��)��i�ћ���v>��*����اL���S.�;�Q�5�v�C��z�c��!�z��w�c�w��Ȟ앓b�wM��N�g� �l_X������Q�R�G�-������fpeS���(7���x=�[=r�^]� �o�EB1L��]|Ȭ�^�' ���g���ih�@_��XDa�&C/[tWEW��oґ$D������`��q�&ϰ�\�)�[�$�U���g�&�F�MZmQ��#��z|^gzf�{�Ѻ�� U�]��
��=�����P�o�����M�2��j�
�LSⳤ��s`�:��,����1�l���o�>R�z���[��ۇ,�[�S*x�Δ*8��2��$��\�opvۯ�Ld,֚[�B�W�y��'�&�����a�+B�\&����H�tn��c"W�4�Z�1ɫX|)r�ɩ���^ehR
��aW��,iI��7������G�j5�Q�J��|���?U��.$�
"->� �i�