XlxV64EB    29ee     c10���X{�u~(�f�Ms�B����^���}z�B���N+�� ���H�����g�a5�L�%uY�~�����	\z,�:u����Y�)c,2F>���[�]|'�:qjR���h�.�N����@��^�l0�^�	%o��J1���)��:+�Z�4s�0o['�u�DsL0<�\D��ڨ,�#�{),���M�TT�xO����j��cl��aΏP��m�TjDGdi���▚��[���T��m��&�N�fX��P&��vP��I�EO�b�(�� ��� �x��but?����9�fnkG�l��Qc�_�T�vJ�LA;]>���ˬ��2@R|�F˭���\6�io`Fu�
��'a+��M�4E�����	��ʐzX�S������+�	�V�"�)��z���k2��s��D�)�慨�3y|�C�݆�ƍJM��IF�Շ�}�D�G5�� ��4M L���
 �,��£����ZY��\P}98$I9u&�S��!JV�\#£� �*��u����)X+��q+�o]��Hy�O�<IB�)�L]�-�f�ϧ<�=w'��\	VPᯕ_"��摚���$;k�ǡ�+J�T�o_yg��2orН���]�!�rq���x9Iv�!{Z5�a�ͳp�uޮ�����0h��]^2��t#�R5t�����E��=�g@)������X���t�.<��7�z�U�%g��Vf��a��1�P|��Dgf��kc�-�;�|��I?�;����{��\TJ��S����َ��&��CPFd�?L��L+��Z�N⦒jm���+��0.�v�3bF^����qr3������v�����^��J�ԼQ+���A5�64~��Z�U�@3�ǥ�lLS5A��`a'l���t�t=1��nA�n��Eo�gs����7G��_��a!���F��f�ر��`Z���`�19�;�ŕ/2T�Ӆٟ�����KD�:�:�-Y�0h�z2�졉��`#̤K�v���Օ9�	?�O�e�T��x���е��<-M�	�v�`a�����S����춍(���vkК#��fkA�(��D�i��t&E�?i����V+���3t�U�p(+U̙3��CN�8����*��m i8K�o���B�m?u��]�@)侩��"o�+=Nx��I���]��C����H~t�W�RfSE�l#�z���D·�R���{a��	F��O���[���!�[�yA�N\k���x�c�N�� c0�N��譡�}AI}�6]�� {�����ܘ;�`_ �Sװ춑�4e�+d�k��}"N�8�3��Rr�^�q�?�W_/�����K��V*����J݅ �s��n��h���4�Nآ~)(ZO�M���ȶ��	�8������|X���KJ��!T���I���_�Xx��&�O3*�}L��~a��&e��l9_/N8H�����u]W�Z�2��.W��h(r2rAƍ�D�-�zn�L,-�� Xh���;]�c�Yiz�Rf����uC���C^�<@[������bb>3�Q�8&��=�����e��ĭ��!=���i������
��r~|��#���)%7PB�}}<A:��%\I���߳a}�XjE<ɬZ[P�pl 9�zv����yk��˖׋�!ؐ���z��4n������B�6���)�x�L���������x�!7q{�x0Q���m�{:eű)b2Qv�ʥ��xU)�&I6'59�=��x:I�2SF'����e�[=v�ؒ�N�q�k��'^~�ܻG�����kpm�o�i����!���Wc����hWW��c$ħ�*}��lMi�i-�@��#U�Z��ԕtL��vg&0(KjZ��/T�w��MO����g�8e�`�4��͉<g+��X���\���Z�o�S)���F$>��~�����cw�tk�=��Ϥe��ڋ;R�����QMx?�=�ZV-l!���0" �~�XԮWF?x��~]��j׳�ˤ|���4��K���q��E�^=
���~���t�n�b��f�(
���{}����0��<Ez�"���s�үK�}�A�X��T���RG�����ռ-�f�6���H�$`�x6�N�v�قT עH\9�	��]L~�tdw(F���uB��Xbl�+~[��ޕ�܀���o'�L�jq-���C��hru8 +��\�%�Q�XaD���N�ϖN+4�Mˆ��1B��tz�4����h;�­Ϟ:n�7_n�Ƽ�m>p�@p-�㎓�2�w�Qx����G:H��-ա9?�ޱe�5��ldm4>7:8��V'C�O"Jq{�_���8��yIzk�1���h��X2�;�0����t��#���W�8o�A�@ښ��U@�u-��Q<XAń��^�����:�6]t���M�H+*�IR���j�eC�N���
�
���Ό"�Zh�YG�pW��w���5�bD+u�-�X���}q���-��0w��>�S\�<�SJZ��j�]�*a�����C/���'*����J��
?9	[iM� ]�!u:�EʹͲ!J�%�{��������?��iG����Pxz��]A���7#u�Gdu'~�%Ptʥ+&xG��
�ݍ 8��;*��"��qt��� ��S6��'hG����1��7d�M~�7i�d��ɾ77�x�v�����<r���#��GC�4���̚�7缺��t�o$^L�ҧ^5���Qn����s0N˲mҪ���gf��L	����������>�%{��&7X@̉�i�
�� �,���#1W�Q����4��vT"F��L��!!�9#��0�*p��~�^_�mR�O2�5n��{b�дvv�\����@�_�u�Y��*�GC�'�Qr�e�������������-B\�Č	5SFZ�5��T2��L�3vC�Zv�}�/$�U�sS��+R����9��K�1g�ˊS�n�B���4�:��h]��E$j�l�!{��W7�2&�I����Ĝ	��C����`�A�Y:�����;��5�<n����x��=�*��7�\&hxx;�-�(�