XlxV64EB    5864    1350t譸~�j�#�)�Fׯ�q�_W<Q�SjnN|l��W�/�W��`�y6|�<�K\2er�9����iυ�8�M�)sף�7'J���iP 
&�Ƭ��GrY�J�çeF0�\Aܦ��b��cx_��U��:�B����~?�!�~����ł񰚐�S�[��$�n��V���,�:	r�G�3m��8W��J�Mp��}��3 nUX�GY��Y������ܐAF*USV>�|��x>�J*�9��abϦ�Bu�nw���$��и��皢;d����&�lϮ�B��A��ռٞ������S0�L#�Gt=����(c�b�Y|��В��ƅ]�༝�Ú�)Nn�@��Y����pC���H�R�Z��4��6�T��R�Ij%se���ۿ��B�-E]���U��W�e$���w� �nρ���u���IkB>�a�-»+���I�o��l�P�����RLS����� ��
���n���'w���d~ӵ3����\��k%���^�M����b�E�ٷN��ґ���]แ������g¸���@ �Q�gy����J��-_��W {O���u��9���@�~�v���A��+Є�>R{�N{��?�Z�,���T*\Yg?]q��\PH:>G8�/�IB�W̓1)A�V�t��[���ԏ���e���<�~� s}Ļ[�,7���yg�
/ 5��6.��� ��j�5#[-c?am¸;'?�ѣ�-N��싚EPLT3v��>nѯY��7�ʓV�Ho�s .p \�N���[�b�3\;NcA>;�RYWϽ�h��,�+X�^��j�x��v e��:�5���"C�yǺ[�-�u{���ǦF�[�f��)CO�;ށ�5�h��R.bs3S���Vw$�6�ϳw?�m�h1���C� \��R����A�M�
o����R�YAx��=^���hIDM&'Ծ$�<�btG�[�!��#0H=;_|�5�.�dE�v��s����>
o3���.���=�E�gx�IF��X4m�+�R��<i�OU?�5}�	��OD�G
zm�>���3�04� �%zϊ�p�6@���R�
�A�>��(e�e�X��D *q�>��1�ThI��jVƞ��*/�±+G%�䡟��1]n����H�'��b��az���~�*��HȍvRN7�4�k}����M�j��h(述�x��J�?;e�D����g��d�.���Ɲ��0��Ye�,8�@ZJ30�o�:lY'���	Hєx�z�N(Tn�|�T�� 5��\��m���sn���������_Gx�[��ͱ��B�o�={������d�5�lQ[�������5X��"��,-g��5��e����pn7DV;�$ѣ��~t.�t�M��/2�V�Q����� 	��ppw��:�w��:sr������~�%A��@�E�*9ɀ=�v��e�^$� ���AT5ߘ���U��-0�S���X��`Yim{Y���"�J䊓�D�Z���R��C7��QG�*��>�$��=�ۧL��[�5)�]g���C��� ˠq>�J>>.CO!3����g�Y�`ũ �����I�R�$�Zvd+?+W�U���^�	��΁w6�4'�A�R�H��7F��D���t��I��T���*���Wm�.짿N$�M}�P�AVl��݂�_��c����������'Ur8�z˄���[�p�W0��]f��S���FV}��	ҵ�o�DŚOŋ����U�ÄE �8~H�3�|�D�A�o�)���uނ7��E����$ﻹ�F=:'g�@+��O�c�)\���VV6PJzҫW10�J�d�:.��/~M�8p�x��4�e�^k�Ɵ˯5�G�����)ũ��_a�+�f��6瀽j�ğ�E�l��d��S�1@�N59���V���)8A��3K~�z��Q�h�4��Kĕ=}{.�<�'K6���&n[���q��Lʥ-����	��%�b�N>n��,��W.�G]i��Z�uQ�`���]��D݀�c����N�8uz��/�*��IA#�WK�4x"ұ2�{�h%J��9�Ѓ��T6Kۼ@T%�u�ps�/�P��r���?���u��B�db
�_�_؎��
���§����J�7|7gWcͤߏy�7�W�&�#�d�
�E��ڢg�K��XڪＢ~TJmA����d ��������gFݛ.F8��Adb��Tm�)S��Q$�A�F�O�X�ܓ_����s�d����#(cs��%{��d�~*Ю��Eb$���W����]?�l�]�z�K%Me��P��5h���x;�4��Dw�&j�wϴQ�k�X���@�M:6�z��F�v���|��0dF�J^��dt��K��U�����*�5���o�'�`�6��aR�Z����k����
j��\��Q�|��(�Q�]�r�����%A�4�0��{JS��m���[K�`0��{�~��i���^���~�����y���%�ϙ�Sȧ��k6�'�O�2M0p�b�f���"���[�E�y�1E�X�B��vE�s�y��2�QM���<w�����Q��T��������kJ��`��oM��̻f,P��N�N>�=p�Ft�PR�{|
jiF2��T��ve񝣔�4�Ɲ���[uV��)\-���7A�+^ր��]_��|�7�ߢKx���2�ax����vj��a�C�:Yd�⍣�A㙐xtݮ����|`�%���*u�y	~%��7�Zt$H#$?W\����u��m��"�ȅ�#B(K~66Ve�[���u��^]����h�?�����N�[�H� �o�c���W�����'�Þ_�9�k��%��&�Cv|ubu�Zg�blHq����Tp�}<���l��(���	�/�L�`0�0�NE��F�"�.%��F�Ea�&��Q��/���G�;��~2���?i��"�J'�V�ȼW�7O�SX7�=�F���;�MU{�\�k�
sf ~T��X��{���%Q{	��Qj�#����R�+PG�]�Q)�E���� �*b���Dʖ��H�O(��l]�
��U�Lh�����:�7s�`����{Rfcڎl;JB�_wNwƶ܀�ha%��E�xp�F1�9��uP��$���.aQADnȆ�q��Wm��E�R��Di��3����cr{��׺�M���A4.]�晋�	'��X�H��z=��H���}����l��rM� %w ���?�ʻ���?�Ȥ
NhQ,��*�$$.����^���2_���|�����"3�h�q����Plf)��y�cZ'��ˣ�����p���"%6�ǮN��A|��R�I�Y��=�{E����L?'r�/�Tm���"]����W;[ݨ&� ��>���ͥ��\�]�Τ��b|����bFh���F4���k��a6�	�r����2�ȣS�����6*AI�6~���������Wg	ȔtB�#�$�)7,�ƅ:4��H��e���恝�o>�\���t�ka�����Wvg��~���l�����~�n,m�	�}�X�P����F�'�Y��hG��&xu�p�'ȫ8�I�|:c`��z��y>��ݞк�nws�ev�����!�A�]>M�a���� :�78�H�9�GU�f����Cõ��*/��oK��x6_�^���t�j��oy�����0YB�(�?}��!x�ݜJ�Jyq{���"�S�T3a-�e05��T�;LV�tZ��ԢR�vK�3h^M��P�3�,�m���:��Y��G�P���-�.�f�����[��yqP(�/���4���E�e�9�1���]j:�s��)��ʗ�]��6�����ŋ� v*n��e���퉃b�X�:�Ef����=���]��2���6��6�G_��ׂ啈�t^��#���K[j�r��L3�2�����"!�*j�˧���o:Uc�[��e�K�Y��a(�3��HMdH���IP��9�\�d��l[#'~Z��o�.�:y, �Z��:5���ŢgFe�튺~l�������[	B��g��V��m�?*�������������̴p|ty�6���Z�(;C
`�R/��J�f�YN��F�j���nr^�+[���J�\�?��G>�^X��k�YI��~�ϴDt稑%��C�D )C�-��O��Q'	n��Oޔ(�C�3����J撣s�l�p�Z~�$R�� ;��3�!oYc�bE͚���A�|�p�����У���X���
�3)��i�������$z�W���c;�z��v:sl�i��Hy�K@����z�Rbŕ;>���0XH
��X4�d?g`Rt0��E�@��q�1���9��?��:E
q&O3b����}����?��z���9
����9=ۂ��������^���[��X��r��S��u���f4���&�%;1��m��N���+
f���{��ia�&���V�L��D�tӡK0I|?%����dH�����S��$���nK�{�?���\�|��$��p�6�M�8�@�O�);�6�X|��<֚����0CNw�a�0�+ww2m}*�\Zwo��(f������fk
��>�Ig��/��@`���
�P�s��3ߌ���c��(k��
������,�8xNJ�+r@�5gP-��M"���6<��CJ~��@_�B��иh�����>����oYط�ozGȍȒ)�D�^ Sk���}�zK}_����a���tH'�B��{d�N�2���"�a��a�