XlxV64EB    23f9     b60�HJ��÷�%.�<h�����I\a���6�QW�w+ 2�LIڿ]φ}�l�b�z9=!L� 7壆������/�Į�k��QS���{�D�{����'v>�Yw���稉��T@F�����fqf��ge���GoZ+	!��Qj˫�ȋ����:��=)�#��$t�"p!��(j��㾻��J��E�m���PF��♷�ۺi��%D`��{F��)�آ�LB��B�ea3Rխ[���#��q')M3��q�[o<��seF�,@b�J��P��~��o��F�}\�@v��ߍ��E2&)�1�d&�q׃]T��f��wm=�bfK]�mQ�.�
���o@e�R�ȅԅf�7	Z�����Ʋ��z�.4¬2��W�| ���j9b&v(���"];"���Z��Z�E�2�K���pZ�O8!?�ּ���* �#lȳ.���E����̺�8�hʕt)P�V舖�����4��gR%a̐���s����9-�x��#=G*?j㗔=����ro_�d����Ӧ��M�0B~���d"s��35 )�z�0t�b�(XL�pg��C�C��`ܑZ�ͽc��ٵM�jQ��۸ڴ���w�}�x�d����7�����|�L�~B�-H&7��~׀��Grh���	='�Z]HP���e�Z������[�+a��
�2�T�||� K �@�Tq���J̜,��X|@�e�ec�P��EZ�7�*���?h�׻u��J��� HB��"lW͕B�~`T;�ǿ7w�4�����{T��.W��Y��#� ɒ�F�K�Y5X���dɸЗ�Yy���N>��6
��W���@	��Q0���1�s�4���$���l�<\�M6��f`��a'�-�4un��^	���z�ϤJk���tWjo*�#Ih�E��|M]�}�dj�/#��s���A,��&�.04o!����G^��;��2����B9�@�u��'B��*�D;�(��������]� o��E��쀗�&?�Z���}��Hj`D2�_ꈡ>/���^�L�v�iY�"�
����֒O\��V� 9�Y�bP`V0h��:1��X��]��^E �z�K}��B�Oi��WEG����y���	�Vm�(�Mc������������ 	�ݜ�ƞ+�q�pv=�!˾�^��6�Ap�C� L�t��`����%ř����d}M���O�j�"ڑ�����k��QwZq3��M�*����y��o�<2.��֏��i�xޖ
R�DU��������ş�4Kzw�6��Vρ%@�q웃nܲ�8T,b�x,���4����~�\㕡��N�+w2߃F]�F��"�?��}�ri-Hx�^!Y���ɴu��ْ{����U��@U#Ke�PX�A�u6.��@��qWv8��O�!2S�sbp��YAl]|��p�r�Q�7�[E���:�l?�-�;�X'�S�[�{X� >w)SX�����r���t�/���!G��-�z#�U͏#��w\�V�!���]PN�N��)H�Ԭ��W���;�a��/@��Q���T2��J��9����)7�)�Q݇�u��o���=���Wdg�J�t�����g��0z��OHQ�qR����f��0>��|���D�n���v�Y��5��t�]��;�s��M٣-�1��Z Q�l��k��zė�-/NGw�b�S�|I�P]�Hx�$�	k�=�̐��8)��8�8HU5G������C�*ޫ����,��1!�@V%:o��{V�C+�o�S�O�b�Y�sZ�C��q*�e��F"vo�3̎!���o��h'6.j[-���s7��
Ń�K{��E:����^�*[��@Waё�Ӊ���V=���n��莎p��3�r���`e��Z�f�*�cN4)��x��R��U}/nH�6��yФ}nܭ�qaqq��ڬ,A���}(���r���z��-V�*D����?�*�ѩ���H�F��'�šW����T��fc��ⶺaiæp�Ȍ���ŇWE.n�`D/�<�,%�EJg �ӭYL�펤]g�uB���A}�W�	��4e��Y�}`KM#�4�D��=�^�L��==k"��Lg�2�xUb=�T6�0 >�Gھ͚�y��,���G�F�Xj��~�l� ������u�H������8K٢�Ϫ��>�΢�����)�
��7pm_����>\��<DK�Z�):�L���H(?*W��$�����$��a����IbF�\���wZ���>鏀��J�LM�ݮ��꒷�Q��ߣG���<#��O� � o�-	;�6� �/�wc�G>T alp�s���vܛ�J0�����6b߅�tg1+�'��,����"⤾ƚ���J���1x��^7'(��Z^y�U���Oqն�^~�RY���7�d�@,$2���?I��;o�Rn�7k�p�ʾ@ׄ�c�q�G��R���7H������
�o���D����"!�	ctOR� .V�k����52�[~��"�X�y&��iq ��;�
,�v��d��=z1ո��u]+:�N��,UgR�C�8ƳP4K�7"iA@9J�b6���4�G��.]E2�CzWp���5͓I�^ba{��Z6�8�4맅��l���{�Pc���6�f?���
X��`����ޕ'���&�1�.�:��eU��	�n�i��'S�0�-�[*����@S'̭5�2��/ �95k�)�u8�b� �6�*��~��J:����3�6^�����Q�()���fZ6�F�mO7͚~*��N�!�+_�'󗦨<�"v�+�27\�փ�ڡ���\e��_�C�i���
0�Î�\�s��
�Q�o�&u'�m�=��