XlxV64EB    25e3     ab0r���zb6��g�OXjgz���F�mj/V����}ޝ���:P'�!.��0I#�03�cQ�~��dm��A�����|�yTnϞ��r��K%��3��fҩ�!]1L�8?U��Ēv�p h����qg����ӈ�BE��X"P�A�8����PX����ְ���PGj_�)�+n(]�D���̱�wYSc�&+l�8���J����ð����v�[��,����㒧�w�H����a9�J�'%�����{b4ƚ��Bh��-��9�� <(�^U@��	�@�K٘�C//����g=�Et��L�Le6#�UZ	J3B9 ��l"	k �L{�T��D�fj��/�*>�	���(p8_��_�jÛR�l�jsӭZ��%�fȦ��X.�A�im�<q�=C��Ӿ}+�`�h��.�儔0�'��?x0-�W�ȅh�Ֆ�����m� �*&�s�_���cHL�J�n�3�չs ������w����$co+oi��K�EI΅*?7��1o_���f��_g!�[���P8\��2.��H������I"�+2�d��:����0�`�r�U�m��C��E�B����+���g�zC�7�l�??��gJ9��o��J�{'�ZD�H��s�q-��u�K���g*��=��>L��eD��
����F����b��6zu�����1ت�[(�ni�f��Nj�F�	�U ���( ��T0����ODvF)����U�ήH�Q�/U8fO����]�|`(�ycU�9���Z�V�9�$�0/2 �l9A �W�Kж"��Q��r܍#�:�N*�s����������6�Bd���D�n�ƍ�)17��ǁ �'B�c��5�8��� .2�O�p6!�ZO"�66x��/>��=`\�S��2��_r��2�f���
'��^�vM46���ۗ-����NE�3�ָ�gf(�o$]�ȭN,C\[�Y�lX�m]Xk�Wާ����ϖ��vW�bN75�~7'{�@,�Y��+5�D���g��`�Sj��l�?�h��:�y�c�
�=��� ��f^}J�l���T	8���x��ct���vg�}|�Nŧ���Ӹ89���u{��x��1SMm®��W-!g�z�'� ����1��<���;a.��+B�?��?9�����u-��vkn s�
*-F� ���%�
��L��w�uatJI��2 t��La|�y��׫H���z�
w���n\�#�%G�閭#L�1"hGsIN�h{�5baG�� v�yR����F�G�6"X�Aq���_F-��B�=�]�W�KIz&gY;ᩉAO�u��
=	����r5��I�o�]��Í��'�9���$�2vRѣJq��R�8_�~� 啈�7���TU��`y�n�6���FYBBy
 ��q9�s��򯺋������!��W%	��|(��)�|&p�8D��A��zF�ɲD�����7F!���[1�C�����$�qj �H	��iѤT�kMbX�I�.�l�N�:+o�34A�ٔX��|���;�����&����������~C������	!fm��3���U���$ut�C6g�E�!	���(mz��\���7GY�_����~u��4�?^N���K��
��w�`]l7#�����Nn���bYN�W)a�ɓP��z��z�uC��530n��˭��z��z\mC+*1|x��l�?8�#���3q7nqN�Ԇ�V_�2�{�>-7"Pԧ�XT����h��sY6�����
�BiPF���	.lTy0s�b�DE
N� ���=yD)�-n���r��7Z��*�F)�>���"����3#��>����n�gY�N�����8F��@%F������q��y��-�\��Ȟ����dz��ٽ�&S�ڶ��]��b9q�r�=��͐���-��b#CX������K�*��^�+�w� L��L>��[�2���0�:��y%۔�<�z���o�W��i%��P�~�68W-"�SvSc����G9��n���G?tsW�F"�=M#Ɋmo&�?�2���k��]$>'i�4� !�����yUTs��6�]4�x�s&{lS|���� l���#�˼sC���o��)���=\�
Q�M�m`�,X#}�a6����z)����b\4	}P�����I:cP��Q����u����h��ּ6٥_���	��͙-��|���˄�I7��ܲd�w�A�&���<ڵ��rt�����`��g��j����>��THR�b�C^��p�r�u�`1EO��)��܎���~�le����+嶖~�QFHi�5�:�,E��L^�M(�=�-C�D ?�zbQ�DH���A�".�y]��� ��W�~���sA�M㚃dC�2�@����m�d.^�2�D�1א4$� i
����>#�zNEg4����W�ø�uP�a4;��11}��(�+l�'`�0�N�36m��L�g
�fl�RH@������WFT�R-��(n��̾Z�,<�^Ka�%6˧#�3$񪌼7Qn�B�y/�E������m_��r��C���m�H�u]4�-�i�ߌ����(����S�ҙ�6P^�<$�^��_Y��+w�ށkI�T�[�yhn6"Q�7��/Sgb�q��}Lƙ����