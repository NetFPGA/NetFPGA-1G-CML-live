XlxV64EB    fa00    2ef0�q�3!��]|buE��<)0d����*$1��fE��G�#
��o�(�X���KԓC~1qN P>��-Шf��0M�ǈ��yG�g(�w���CC�V{�Z>�G�����P��om��\�d��LEn8��d&!>[���n��U��̷a��U��pְC�.p�u�0�|�XEύǼn���g�YN�髣Yq����BXxSkj�#�� ^9�����wgy�;�	��e�`9�̇�����pJ'�m�mr�!��5��2,���ov�P����{M+��m�1�%p��t��} �O�q�߹�oJzL!�_��I*`2bR�Tt�%j$o����G�W'�WeF٬���%�,��Z�Kr�F="J�:��
�i���;ߺ�x�}L�U�|L�l*������#mu/�*޻��#^C1I<�j�Y~fG�����L��1�v�+}�8E�g�����wN����=�O��u��y�պCPB
���4Lĥ4�hO��YCj_�(qK��$��6Pi>$��TР��ڮ�RyA@�4\Xdn�������+���[m���>[��:�������ϧ�y8f�q��{�E����m0�Xo��-���;��/��^U!����E�Y���y��\���$X v��2˃k�c�%�zw���&�R�E�dݎ��8�kk�)�[�߼��;�kK�u��)�h_m�ԅ� ���n�iaȇ+W�16�|QS_5Ȉ[��DE�������R�!�Y�`6�g�����x��2!���Ǉ�G�l⡅���Kۘ�x��-/t�`#���D�A��Z>#i�ةIU6$*����U��>|b�|#	>o-�vx2��@��f����dZva|���r�ޡ�K�Aq4��$�?�|���$5R7�	�
ps߷8��Y�;^8�r6���`�[m@�BԳB"_}������K-�X�`:8��;oI�	<���4�6uL�U���>~n}Q"�֯Ѻ�@��:HT�	�K������+[s��kgҌ3ͷ�&�L����I�eR�v���^�	yD�����Z�^ms��{�'�}���%W&��V3����S�&�Ȭ|�i�C�}��Ai�X���kV�d$�H6�V�QlK7S���fk7��:a�� �h���D��Fg�
����bi�|An��8o]�D�'n�F�5+�O�@�N���mQN�cc0)�-]�ۂt��Z����'��x5/�e)S��J�+�co�����z$��l������1Tڑϳ&�Ǽ	#�֥��[�l�Y6���w�D
�@+�fS�*��K�9F7W�� ,�-C!�/�-z��u��`��/����1��xKrϪ��⮳3ŷұ���̵�H�R�ђ~�v���W��UGv0���>KjFY0�:�� }nE�7��G;|.��i�-���2�����;��Vf��P!!�7���!�K�M�n�L"ʈ'Mt���m	�L�jV�|O��
n�x�졥}\�m����w¯�C��ps9�/�/��J��ې���Z=���e��n��l"[�oA�g8��A���R҃����d��wb�Xp_��dА��q�a۽7�9�;�n��������*R�`(�_jp���;h�t��9�ka��/J�p<lQ��åYKE�й-#3+��>=�&K��睇~���]4aƜh��!*�5S,rMcޏ�Q�%�C��w`e�6"� NOcKMj_����V˥P��c/������"){�8��)o�+���l������W�����=�g�z��7o=�0�-�= 0�
�k'���k���i-�dP`�9 [�&ß�!���������Yc���Q�%��AX���/����Q�,!��]8[U|�Jڝ�+���S�d�6N^٬���2t]��%=O���>�a�.e-��׍a$q�x������_����]��Q��K�]�/�?+#D'mO��t�#������方��K����\|.��o���F�A%B��j�2�53���Vi�0���mNz늽W?	Fm�^���|���6v�ƪJL9��:�Yc�=�r��+,�����t��gT��Ó
�z��@I�Z`��5�v��1_4�d�/egT��q��sCR_�gS3�#�������پ��C S��v.0�,EC��p�������-�HW�Q3U�|��:\�9��⫄��x�\$������n��qL?���W
8��=˲ۋ��G,Ì&F��5D����&�ۃ�~��@���Wo�ryh>Q�P�	g�0�_c�$ĆrCަ�ԃ�ǭ�*����[�y�?�n͑nx�ǹ"�:�'�|��s\�rw*�Aq�w��Ǜ�tN��G�m,=ܜ��T�����k�{�j�À��AQ�q�w��R��T.+\,��0��c���zZ��u�U�Q�f�37�}sBX!�`��ص��� ��L��j�M���2:��Jv�eٺ3��򹦞���iӯ�t���M� /� #���j��Z��g�-2g���6{�Ԟ)��p΂���<��+���<�R�q�)�y�G�� �o�r}��;v���7�����h�Y�x��a�j<ܚ�q�y�3�d@��3ȯh�l�R�DKK�v�]qד)/�?hs6}��j3�(�G&0���	���OKJ�$n��d�U�����I��"�OX�������YW�(�"�������Z�83�^G��˽g�4�'ZSl�˳S�~��׵eUXL����J�Xs��ѩ�.�F���w��p��6���F9���"ݳē���
��p+�
�.�E:�Ʊ��#��W�q�E/A��'���`=(O8=��]�_�S�t�`�r��6�����K W&	��f�f�
Q4Q�s�Ti��ta�+�A�g�X �,N��y�1���Y�!�
�&Ē�W`����vz2����ɺv��!0��ʰ��z�|��u-�;4�Aƃ_&�����DEjF���Ofok���2F�@���V�ѳ#�1\�WT�1܊q-�̹|pަhQG	�@wc��C��wcำ�h<a���>�~�+V���i�扒E�����Y�s]B *D�p���j�)�${�T���⸃��$�~1"8O'�;J��G[wv�x��fP��]јp�"�p��1RSw�W/������2��1ɳݭ�i9�`Ò�|f���+4׮mG{�-z b"�g\���H3ĜH�����=e�5�������L�,<J��J�9�6�F�iz@3�%7���ڹ��=�dI��7ZF���R��m'n���ٞQ�@���5XJ��K7����4'�X0<��`�Dc 8�ñV��j(.
'a�WH\)�d�h��,d�Ш� (�ie[��t�6|m�n=u���q.qk"�a#��* �x$g̤���@��\�q��TvJ� qQ�).��:�/Guc=���]tK?&_�Zyt�w�=QY��D�n{7�Z��lp�"�	d�y>�������W ������q��_�ؠ��_����شv#������D%_)�fe����֘�|���@T�t�ح�Jvk�	��������G��yh^���<QW��DuZ7Y�x.Xu���/�bQ�n��Q�B��{vmO�M�W���,t.�.���d�m��u��ӅĴ驼��֑w�)������΄ Ŭ��x�2 U�a,|X���Q��iH+��c������u�-J�S�28�/n�LD.����ˆ�I���1�8BLX��1𱷐ag@l�5��8� �%�G�������!��"��}�
�H^ζ��n3��B��Ldui[XO���q���)"Ew��2��[ӥ<P,r�c���ۨ����}W��K��	�P-��8��E���L�0\@��Z�%��@X�����x��]-�Zie��QU�[Z��Z���Bߝy|wV��Q�s���[����Y�kgT����Ú6_�1���yʠ���t�-�]G�����q?:���n�g3�[�� �BV������6s���f0�핻E�TS@����&����)@/����AR�[�����>�.��G#�����-���͍V��+���k+�]����,{J|����k�r����
<v*����0��H�wD� ��j	����x�.�����:�G@��=H�γ�L#d�w�v#������"&�c^�рHv�-�y�Ԧ�z�G��e6�@΀��hy�pX�N�W�ج��sIC0��f&l�5���7]{��#�1�|���k��f��m�t��!q��\# ךԎ(�Y^���~�����Y�Zm9��pD�)��t��@D]GFt�c�yZ�Q��U���q`"�4��mi'�n�n��^=�|$GD2�Þ?gnm��3�SQcp�g�6:m�mZU����J�����O�WL�p�Q�`�b��P���:>��b�����ע���p������ƫwKe�7�7��
��Q��$��+���8]��A�{J���P�d�C�e�{;[������|�7�W�{i��]�Uc*�a�7��6wv�"�\H���(f.���c��BQ����]uu���S�N-�..Fg�9���<����$�$�>�벸��j�Xߵ�a���J5o��4��2�,\��5�7�#�u&7�Q�W����K�^�w�1���Q>(�o�d�ۼP�=>�H"d���>05e�4��1��[ܵU�υ�m�Vi^�.A�0⟛.1��|EQ�Mm����=H�N[t�-��v/&�r=�է�����l]��F?��.( �@~��9X�m�o��b���2��Z��e�R_);mE�y��:%��&9w�t�? C�~+a���]���.o8;,�?��~��]�������U\�����Fa�Ɯʗ�� z���P�cp8�H$0�d�[���c��7)�MK����)MJ]v�-E�"zRkW1�V�س�Fx 2+p�bb�py�����Y���4<+��=�{�#/���������sDo�_��!����5��Gށ�2��}-1t���` 	���	�;��n�3\�g�]�L�|�O��HM�O��f͸i ��6���IF�ttI��c�Тh�L4S!�A
oPuQY�j����������_o�?.����YΧ�3"���j��y�S���RM\��7|�O�L�*8`w!�4���̀�_�ʦ)�}̣�=j������`4n0��Hk]�$Pȯ@�� �11�7? j<�w�q\�`b���S��'���������F>N.0e1�Xԑ�u�F�l'".���R��Oq��PЃY��#�����s"��Dۋ4�}JĖj��
pYS� �=�^3�g��'�れ$e~ħ��ZX͜���=s.R}/	�md� ᣸�b�-ǸE��(V��[�� ǁdo�2��v�L5x�����!=��!~��.�ڰi�l��՗�C� �K<-l��$�+"*��g�j��#�%9�x)��ز��7����.���|�ڙW���ѭ��+XS8��m��8E}À��m�A$2�_�]�`g>)�X$��vħw!�*��\�v��{�O%W!~�'�o�p�������z�y�)���qʪ�7
笩� �8���^�`���.�C���{�����&i&��GD{Ϧ��� ��=}�P��=F�?�;�&�uƅ!��Q����Q㳗���:��؎��̖/�Z3t�ƿ:���I'Zw��G%9�B�)>e*����,?�H�]!�	�u�ϗ(�*+g|�ͭ"k��Aɲ��珄�n�҃U"w���xʽ^oH1���L���Tr9Vd|8|?o��#֜�W�+����L>4�+�	�}�f4�i�����B� ��;>]�>�|��?�,��(��/�]tx��"U�f����ḿ�Ë�/��`�9�/�*�G��ʖ�zK	P��iѴ��9��D=m�)�S*�"�8R
��H��n���Ы�h�-�
��{x�QY����O1�*��9*e�*6[�2�3��������]�����^k�q���IM��vz��� ��fXEt�1&�>������o��n83�z[��ʇ��-sN��̄�h!@Z��F��4�����zw"�K_6J|9q�Ec��w�>���麡���Up�a�V{��gm�<���je��T5ā���\(��5,A��À+=G�G*�1U'��ջi��|���KM,NKS����D�z�z�6[��>Wܳ��Ly��o �*m�S��uTO�Q�s۝�O�xl���r��2-�����w�	���\ �W�8Pu��������z�r">ͯ7m��s�z�b��Q�foR��2�H9ץ�R����^YG�`���̺'#Q`�9�]6z�L,����<��E��h�bB j5�BC�5��c�Z�D�DZ��ԇjZ��/4J�ST����;�_ض~4o
-�Ύ�8��8cD7�3�Z��w}D���~��J���zON�@�����El��,-=(��m\�r�U�0�H
zMYT�a�y ��wlV9��z�YPvT��k��3��S{�u��82�錶$؁e�&5�IPyB���V�R �3I � Ǌ��w��
3��<�mi~Ө�?~.����3[G����}�'��pW>��_P��EU�+��^+9����BCZ����h칏���]I���@-涘oe�
Zzt��E���y�e����mf����_���Ѷ=ǂ��RDG8�#ӉRW�9�Ч�����j�����>��ŧ>"["ў�a���S֑ɗb.S�-� ^r�|%��Q�
�Kk̹����j�I��n�]BT�)c8E(R��tg֒~��1�*�@.R���&wo��>� rwl�}��z����]�!��@A�B�=9r�u�>�����XT�.�O͈��z0I�~"[�����Ȣ�b?�k
� i|� &ẛ�|ș_O�өB�� ��.��!�f��/�O�0�Bݒ��� �O���:Q4*�}�`��i�����F��i���=���=�Ƨc�Z����k���X��ԗRy�b͟�1{v=~i�DhF�졄&��#Eڱ��%?����v�������4$�VB��c�\�	��A�+�Ơ���XLI{�{qƘV�i>��_��h�=t�ˮ�{�� a�?�=�8���I�֋�譣>�l�` �q+���A��a�O� 9��� )B���͍B	=^Y�،����8�������
 ��c�F2�Z72]��MŜ��ZO n VN����
���z��'�j�L-W��[�郸/z�#�/5�ϰ8XS c�s,d���&P�`S�PPԃ����U+�v~�fŲ�m�}���"de-Fp��N�����koMa�nt�>ke��Q��ŵ%3r�����l��08�I��e�o�<�]����b�ᄽYr���.�v��� \0�YN���'�;��N�A�	�p*�D��,�!k`��>bq�
�~�k��aZ@?.s��Ep��_�'z�etO#�\���Q�M���FּT�W���� ʃ�M����I�l}́��IO(��X�+�A�^�ᮯ��VI��@�r�1�H�"�#a�|e`�6���\�'�q?��)ζ��.�9I����J��`�Ɍ��	�|�8�`��ЀA�c;�J5p��G�N�U��vV�&��o.�ȟ�պ��i�2\��ɐא�����_E�qi��)p�8���B>�%��/^���!/=C��٧�@sX�0ѷ��h�WJR���$�+�P�x릡)W���e��-5'�㑏���;�~6�D���'��j���8aЉKz=�,�s��X;&^����~����0�Юϰ+��rt��h�;��5͘�F����f57@�h�qY���{e�tp�t�����Q�@$�-&��^��
�峁>trY��崠�R���_����ߤ����dŦ�{���,>T�]�OB��u�wx(��kL���S�Q�:$�8��3>�)��d��u�
�%h�'A�c�����->����:e��L��x��:���ݜ�ÀD���)4:Y J�j㟢P�����:�I���6���%�L�c^ ��Y�&��qt�S쭿�Q��������F����fh���
$a�뤗M�����i��<�@�?T�2���+z�1��H�N�8����@ҙ&�0V6�N|-�F�iN�ڳ`�v�\g<�(���j.e�^Q��z�GR܄����1\Zu2��c�Ꮒ�A�;���z|5�5I�t�!�ytG���R8��M%�,�M��G�E�'���r�9��k�!�)�^��M|�ٮl�E����5�g(��G�.G��C^���<TPeg�^G�r�C����p\eK&+��<����u��xf,1�z�f����`}�l���f�?X�N����S]�$ㆍ�J����XR�H ��*�'��6b�Qu�3 �-dH}��(�gi$fq��]R����ɒ��MVMv�YK�t u�eXfm����Q<]�?���o#.��|Η �Cq\,i�G�W��ؘ��I��i-����#�B|�hx� R���ǷS�e�NKZ!=�%��6��K�'��ƖE'�i�*z�0m�YZ��c`��hC�R��]��j8#��1-��ː3�I�j�m��}ٯ]L��rX�Z����I�.�0�+��`�H��S��_����<Uw��((�����g[#u�[؉'28��PV�5�qc�9f�!?.�^�P�n�6�w�Q� �˛�� K�a�����9�/�%�y<�Z�4[�B�{4�NK�)@��݈�Y����$�n+�A��u_+,��F�&TBWF'�����v�W�\s�KB�L��*9�����g6˳-S������be,ԩ!��SL�500R%ܱ@����$��a^����+�1���ͼi$֔	U���7���W�N!�N��g����(5	���I[��o�+���B4���~.C�s���IJ�,(���H�(U�myT鬪](i����J$��e��,n0�j����_o��5^.��a�o�SA����X���WP�<n�\����O�LzWJ Q��K>�47�.$��^װ��
���igB�һ�W��w!��N����K�燺��p�Ӛ���`A`�ۑ��~�h�����@��vw����g����7=�Y8�����]Å�3���B=N�6�/�ᚢ�f��{�2M3rN4�P�
���Lq=_�����mG��+B� S���P;Ѡ�-̸��K�N��y��~��|<�Wߧ� 
@�U������s�i�C1��{z��8h8~�j'AC�Kr%$��dLr�	���!SKm�I��~��$�mH@[r�6eW���T���Ә���-:��%�<���N�`�)9����ͳ���xEۛ����&���48z����2W��Y\�$�V}Ŋ�/�>t-<'�d�ܪ�[~��wݣ]���35G����\_ 	�\��Q!�+7B(�f ؇P�Tu�]�f7�<d�_���38�L��Z��g��C����E��a%R�`��������/{�P��K�x;�����
n�l���������WN�O'/�0��� N�bu><�߷� �fA)O����0�f	�h����}W). � �G�K��[�����!�v�X���'�+�k����4��"�_�W&���$���IR��W>��_��A�\�o�gFӻ��J�)�cӌ�>���	[�]Bo��b[W+GO�e���Μw��,Yo({�@�'|zڴ���u;87]GQ�+;(�4Q�;! J)��)S7.�
񗧫�e�_�+��o䴂I`�ı���+2������� ?�f� e����	Oξ�*4V>���)���6��z1y����]�dt��W
���R�!Ԡ���^	�8n���@�p�d6X�&d\�v�X*�BE���в�ժ�Q`�z����5l��`�U���iE�f�8�.�D��Ǆߗ�@>-��K�q�(��o�b��Y-u7F��,�����b��>�摭B$S�]K�"_D�(�Iq���NZ�蝦V�{D�%zglX��>�Y���F���A���j�?-g�a��t#9�K���	���2�\/0�ǖ '�x�������I�����2���OG<�q���bW �I��{�N��d=d_���kz�|�ݘUQQ����҇D�Y��	�t��Q�\lǒ�i9@�+���~uԋ2#�(X��������}A��%�9��	M�6��1+�]�̽�>�W��p��	�$4�r�m�v�M��D<�>�A\l�x��V��3v$�����/�T�)�U�d2��s�����`]��`S���Y�y�p��+) Z���a�`��:XC�L�¤�[�J�e��D�m� ��f���j`�5<���1�`O_��}c���Y�aam&h�u-��܄O4,I*�o��f%��>�M��"�2�(��u�F<��G��<.���ؑ�^��z�9������V�!���	xt�y2X	QE��;R��e�R�LeQ��uӠ#�[�ࡂ�3��CR���;c-�֗iHYw��I��I��Ro+``��>����Us���_	j%��eySf�
)����d9�QV!kg�O7 iϫ]�dd7�2�  T;�7��@l�tS���f��
r�����T�-�<�5,T{'�s��B�q��l��D�����u�$��k���痒����.��K0��* �J�B�A��e�X �xd�P��i�ye!���϶�ۇ�w���1�N�^E����h�����@�I��ʻ[ӓ���/p��� rMC�&m��ՏҾ}3����]AGb��sw�w���W7%�S0\��"�[��=��)�	��
�<�;K��,#rÄ�@ݯ�߂F,��/6d����c���+k?XTwҽ�?����!(]�Y	��2g��K���'�#��}�$��=����+X.ɺ3�n%���{�ȗ�9Ȅ�f|�X����)�UDS��g��o����-'Ŷ��a��)-٥7�)�JU��� ������5)0�~���n\tDe��i���SMy(P�T��m}P|<��}�`O+�� �y�mLK��r6fy�ǄJ�ú��IjpA� Q$�\�.�����|���6�n�e��_��y����&JY&'0LzT�L����B�6�L���֠��2�'�/r�'7?�vG��#���o��Bw^V��Pm{�Ѷck�)�w���U2�Ӵ��acm�떘�B����b��A���f	IE�E���Z�;[��eL:��T\8�ι�>��5��r�+>-\�z�,�!@p�grl���ʡ�_Mi�=�|2��F&8��F5��̅�H �rd����(��x1<@���=E� l�/�S)H���[ӭY���.d�gC]z�z�z�n��}T��Ĉ�[`��]�$�,ER�-Eܠt�\�i!Ķ�f\۝�}��������C��_66��¬��M�"7��u,Lx���A�Ս*f��R�/��U�z���U����`N[�HO��I�	�uc����K��ء�FI�a��1���OMV�����v��o��0�v�����n�5�sHo���}V�C�B*�������걤��pU�}d^������J���f�w�	�S�r����g�`!�&P�\�����CB���d���	X=^g�NrZj�'B��iOw�ʖ�D�'�<IV	m|L�ҾX�勈QNz�#���� �@2PkY��QX�ǻ�}#y z��Uݖ��"_���Z dH�}�"���ٌ�Z+��[8&�y��I�i�]����z��fS|�n�Cz;!��B�o�N����cXlxV64EB    fa00    2be0�eqh�r�A�H����Q�`)�Ϧ�Q���E�T�|�Fs��B���;�.2�A��쌞�(�#��)ܐ�� �ьȁD&Ɍr"�n��bHZ�E�O��Þg��PoKH=�`�;��AP��y�~��0��d�lG�/:Y�;��#�[b֑S�H�(e�?S5�;Wr�_�oD�0��������X�ە���?��u.�cX af�HZtq
��@�F`��M0V';l\��Rk���D���![�ȇ�b4��K�tsb�l�B����mgC����D�����끵�5޸�&�TC���lZTȣ�w=av$q�޹H��`E$��lp3��qx-:���4�S��D��L�y.�0Tശ*��v#63�On��E">�B`������Cg�s>���9B�e��+����7eb�	�0.���w֬�,ԩ�Ǻe\bt��4������˪�nEu̷��3���2ޣz	�[��Lޯq��p�#ӫt�yE{��hh9�ƚὶ�)������l�[$L �_n)]�O�� �Xͣ�'���".���sCD$Y�7�P�n��&o�	cb�P�`
����;Ī>�2���R��^!��o2ˍq��(\I2�KO�$K�$�#��[����^BL��۾$؃Q�����v�w�#oeR�����5A��w�R�U5�F�q���"[����or՗�WP7"����~��>���������:g<�	���M�i��U2�l�
q�b�T�!:��6���Z*���~��3Q�`:�$�s��r'L��/ܓ� ���;ã����.5l��I�{T�_L��:��1s�W��Ba�-�STՅj{�桜Uf�����$��()T���
vj� ���NA��J�Ap8�o$�h�ރ΄=2.I8�'�9�!V� �8�h_��6*��m�����8��:1�����X�ꙑ�
v�<B�׊��d�f��!�#y��N��'�ٕ�C�q�pV��8f�ׅ�{���q4��.n�c+�ϲ�R�Tܥ��G�DCg�Y��� ��F~��3ɟ����A��W���|��W�_��)T�*�D��|�mx�������r�@�)���J��*��N���N�kE��#v���?�B~����Ъ�Ao�%zRA�/�	lw�y6l�\�t����U�F�7�<��D���gS�o�/��'��x\%cn��-�Z
F����Op'�zi�u����&嵡V�����Sp��ڹ�q����nk�"���^����9.��xYba��)KW��~Ϻ���3��J ���B0�P�sŁ��/,�<�TT��"���C^�3�º��o��5�K}�L���$�����9��NM���m�lb�"���S���f�Ȟ1g2��1g���<���f!�S�mbh(���wo��F���!^&��\%P�����S��K��Ϣ�>����
�7�U}�N>G��D�{�B�lӯ�T��`\�s�N�-O�e#�a�S���E��4�,�X �F�I�����2���=�gO"���2���T�L0�xʐ����~x������M�k�9bC�L,��IH���S�T��D=Ɇ;X熗OT��ю�/S�A��F㶟�("�L#ʝٻ�C��f��_���;Trb5�!�
��9� s$����J�7h�Ӭ�|���9�b�ݚ
����)T�[�z�:R;<!�U�������^����ΈP��W�xK�~}��j�w�8�<z��F�}��jc�����y`�ЃCYR�g/����'����h�8���;��Y��/c�S�VqN�d��}rN�\�ܿW 8$�N\~\�{�nv���R�uF���Gd�Ό7��:q���� ���g�'� �3]@��^�^f���S�d���S\�ȿo.�oILxK�t~:���a�i�	5!s�s�
���^:6�8t����[ qS]z�Ӳ~0���5�=���-x;˥)Aަ�y�o��1y�X�F|om�iŢ�;��X�r����2K�����D �/��H���&K �b�x��+�Q�;}�[_� ����f�b� �^����/�p��7��o:˪d�:rH�:����s�;*+�?��tC����k�œw�6�	����U{�Ƥ�1m���u�^]�@C�swbWa+����$��p_�5���Y������?�2��Y��p�N�z��H��t���׫TG?�3�ou�T��EM��PV3|��No��W.nL�q�<OܯE���:t��d�|�2�/��P�mt�1r�QnXd�*nq���N�����>N������;h�j���n��gᎄ�Su�C�����i����7�ֈĹ��=�����1V�����d� 7+�u"P|e;K�0��*�X�;��4�ǿU�*M�1����F�~y��zo1��g�e�r���byh��le��B���R����V�c� �g��Vl��i�q���,bژ���;�2��NLf�#�P��X����v�Nƒ�U�S���?P���;���v��µ\��yC+Y�T4e�i �>⹇$ׅ֖*lޫ\i"ʧw��<ۘ?��u�r��Z\�U� ���~X�b���I�W%���a�Ӌ*��eF ��6�G��m+��>s��Й�}� �Ip�8��<��W�Y&Z-S�W�� ��r5���h��a���nr�B��5���9b�����0����*6,V3�dʆyo�Ԝ�:U7[Ł�k5g1�-���c��Qx�pb�h�`�ՎAv�aà��uV�_Blk�9QE�o��5��	v�4�
1�x����J'�9D�o�j�LA`��7_Ц%>4����>��7�L����k`뮖�lil�P�9�j[ב�v��QY��=U;ޒ�Y{�������~s/����lL ��-���z�d��V����J�z��c�C	pߋ7�-z����"A{I���^��)����'�5Z~L�Uh�
4��0ʤ/�]�؈�E�MNn]jniKT0��"l�My�A�<��=���;
����O�l���jD>0�4 =�5�Z���UYb ��nZ���S���2W�>6��#C=�O�3WK��r��N�1b`8��>øٔ��>>��M���8Q Ċ\9���g:��.Oّ��g0x�͘��vQ������{ݛ>�+��w��2,`
����i8�HD����U�. �J�6kҞQOm-��Y��˹�=���Cz�U�f%Ԏ������.;�Oˎ�"�\���P���D�E�J�K���w�{7��T��*U��8�yjFN�m�!(d��|�l-ơ�	�_)�8�&d�]7Tϲ��w�}¿F�{�:�[�ĪZϑ��6ȿ��]?��w���HÄ��ٚ��8.o����1���Iϑ=د��[[b�_ń�&S��<B��D�����m�$�����aL�CY�m@2������*x��&d�8��Z��%r{cG�i`k���Frv8�-�����,���e���8��~j�-+��鴲��y� �g#c_�^��"�D�8~j~uz��'�"ded�������G{�8������G\yz!m�(���;J��?Ҿ7K�]zc5�؉�=�ʰ��<��LY��֖m��H,�p#��k����nj���j�J�H�L�%������j��w|���`�}=G��&fd7N���AYI����.E�x�F��&�� :�NL�6 �S��ݍ�Ȯ���WoD����0��3Z��ey\j��R�����X�Y~��vGa��>2��jP<����UY�Z�\|i��ʥ���u>��v�.I&����V�ԡ��jZ���d&�c�ɨU������]���%����]-�p�v�=�Q��aцt[���!��M�'�\KL�E�͑�����A��ີ^L�� �EFxw��0��;TU����#�0E@v�Ln�W2�/j���ɫ�u��5���_*��}�z�Ԗ;$��aC���P��F�^�� ��)3��E�/�|b��k� ��S`���	�]���b0Gȓ�I���*��N�}.��a�����=
 }$
�p���-���:d�/��AD}�D9�qu�kMڕ�p�܃����������x��p��i�a�[���Z�E_���"S��O�*���M,�B�r�l��C9��ʆd��1�
<��]�x�Q@9�a�k$ޑ���e��|kҩmO2�����>�����M�����?���J�1'd��I�=��-�I�~y�<6�f��R���L���Wg<��B'97p������	3�����|����I2~��>̛E�8��۫��K+K~�h�5��񪹚ѽ�.��V(�'!��2�=�~R��'yL�3Z�Ӧ��M]��(�V):�^O�!.g�%��5�N��Ƽ�*�1�I?��D��}+�8=d6���qZ�"YR��g����ox�/�,Y��g&xɻ)��4r����p����?�ت����A�Q�+vQNb��D��i��W�G��uȁQ|���[��SΒ
�n:�ņ|c��~��E���ZO\�!n��˻&����W�3'�6�9*JWÑ��5��Ʀ���dG���QV�;�;e���8-�YoT���ZlTi�F�+��7��ԩ}�h��T�q��_�m8?0�H!�U.�p��L&�P|{8��V��27��
�tM��y������2�A&(��%]�vP�7@�p��{K,�C��S9�|�?�c�*� R(k�IS��A����������_0�A-V��Q���t��[�@�>x�2�CU�4
��C�k�cv\&�e�d%�חE�ˇ�k�'=���(��FM�0z��Ky��1����,�S��� 8�Y&���y�����݋�2l�x��F��!�$:�s]_��dl���)М?��(7a_2�>�{��,��G��u�
�ϑ�M�׈e?
.���_"��?uH���P�y�Gy��̗��3��t��^��[ӲF��m�u B+qy&���9%��\������:��e2<7 �4b�ް���A�vW���F�K_ZD�����p:�r���.2\�x�xBL�53�%��Z�4���h�D��+2a@�[f��5#\�{�2�),�9�x���V�m4&��_���� B��¾�O��L�2�i	"�����'o��1Y^/y�ըR�-��)�����Y>��,'c7Ճ���E�Y�f��cTXe(UsHpZ�`�^��@�s�*ov��`�׈��N��E��l�r�jQK�0�|:�`$�����]����U���4c��'-�6��9C�ܕ7�^E�O����i����K�bv�u_ms,��Ǧ���W�@_�Sڮ��;q�����z�����)��ʕ���ws�$UQ�	/�4�:5p7v�;��"��W7d�Dx>3���I�(�� 
�44��	��^T��j��=ݤP�|���P[f�o�/��O��Uj���&�z�'wy9�+?��@h��Λ���T`���,�M*Wi�-f�n�c�_�y�2c���g��v�Z�Q�u~�X`����Uܯ�o!���H�ł|���QRT�E'��e�| ig,8%�J�j5r}{���Sz�?�k��m��l��fب9��Lv��Z��N�C��t�ܿ�&:�k�`h5ؾl�se�T��0r�x�d�o��\'��lvHkL��b2�}�{!Z�=��(�cy��nHz�QF��G��K�(�������n��}K����
��t����At��|V�
>l��7ܺ6%|�F�^*��J\pR��2�,�=@�����	<ގA�2
�6�h��%l��FȲ����n�!�S���r)�������-�f��-��F�"G�X�e����h s�Q�y/��í��ё���bd��Mn�%�D�Q�ͨ���?�7���!o9� �ܐq���#�ᶘ�k"J���cc\��L��ݙ@�Fp�·!��mn8�AOix��၇�j���ߐ1*=��~�u�]�FK6i)��c��WcX�����L�V�HQ͵��\��/�u���D���PP�s�09�FsG{�]��W�p߬T{4kg���!����$P�����2*i���� �Dc8f>7XƆK�ec,x�暺K���������~D��(y�Yڬ� ����sȅ�1��?�2��� ?a��*uA'�8. 0rl�J�(��������GYz�[���sa5�b�d�dN�M�v���)�� NA�ͣ�w/P0���e����%"o���X_,v�3|n��'ȑ��Y��f,S��g�xG ����|��	�no5n9�XX]��s7�H;���G��	����������a�/��p,V�����Ie���R2�U#�1��ޝՒ�ۣ�1q��w'W�|5{�l�Æ44|�A�U�����s�7���]|�|���Yj��Ώ B~�M���<n6���fR�)�;�@�D��+��20*�*���c��� �%���=r�Eυ��A_�3t��*�j�H���S��YG�bR������X��;)+�Ս������=��<��J|�i�am������]c��#I��z�yO;ژw�,nA���NN^�^�3~��
���i�"K�7�:�"���U����Nj�0�My�Q��.M�]��w��/�����������)A�\������Dޚ���FZ�W��)�q�v8YVGD��8�7UP����Vypd�����\L�ԽT̲͡�~��Ak��R�{p�j�7P�㽝��7�W��&��ғ���<��ei<� �Vޝ;b�{�t�nw�9�	g����܃��ȟ�㳓�`NH4�����2[�Ӿ�N p^L��iz��[&�B{{|#*n��BȒ�j���5<.���Ċ���K�:������/o�'��
?�{T���eq��/���uqoR��E���n�b]��׽ö,��(�:Hrm5�$��f����( ����9;� s�������A�q:qM^X�"o],�x8)��c8D%@��pF��LI�_f�B�	)�U�j
�����N�Z�o������J�E����/,���&��*�I��w}��S�u�T�{K)>�v�<g�Wa����ٚU�?o�7+,��oI���j�`x�]C�/�^gG��ɚY=d�&�z�H��� T�p��Uuc��G�-�'V�ge���r�in�����h�k:������@�
9=u�y������)U/K>+^\D�f����\J����ߧ��p�ghW�������S�2Gq�jc��iS�x�bR�|�Q��L�\��W�>1%%�Y�w	�5���~�E�`K7�W�AZ����J�l�����U����h��ᆻ�P���I�׆55�Uy���܃�m��L�:�F�R5�=϶u���m���ɺ�������; ��h����mYF�нjΨ�68ˍgr�j�B(˰�/��=Ry�/��ڞ�f��/ZRwUH�r6,7��@xn���}��Z+B�Um�^&;}��*���p1U���\i�ħ���(R��&hj��K�jf$Og���sH�!QU��:�q?p���,�.6p7�"2))��(���w�߾��L(	�r�|��i�З�-n$((��=��e�Z!bn
�����ܪ�l��,����gM�	���ﻯ
��F��{�@��}�-W��APsW��b�l��1��2�[�R�H�hZ���@>���T�~G9��9��N���<�t�=�P+�L3��u�`���e���N�d��ӗg=zy/E��F-���l�{P�_
^���`9�+@�^%�sNG8>xE���)��L=�fΆ��'b�4\q[�ˉ�	�#̋k����A�������ΰ�WuipZMټ����E�iI�ɪ��Z�u�)�#�9�1L��,���hv��_���PqcŴ��f-syLo�*8R��1�]�l�X�^��#��<ԋZ�gS՗��#" q��0�Y2ϕ�U˧c�{z>z�Oi�� m��,���X�N�,Z�N��N�X/�$�u�������:����qW�-�mی F���ȉ��#y�MK���(��`�3��""1J�Pfh�e]�Q��w}&��F|�h!��x�9���ƪ�0��o�'E�C��E�|xp\a0�x	�$�G�-Y����c=U[�J`�i��X�9�BwHb]&ƚぃ�C����IӞ(����Շ���
��iC,܆,�FM;¯��p����RV�g�>�o�����n5�����-g�!��ue�a�L7�첕ALm6���VB�*hb�p���0��'��lqaKxyv>�It�s��H��)��BŖ���($��uưr4SlΑ�L��*�g�ld\!%�wJ��\�z�
�!u{������{'�7�C��Ia��P����a%��+P*��(&�麉O#=�^�g��A S���}[�u��-e[e�ۨ����
-,�)Xʏ�Q����K���Ȩ
�w�c���MπV @7��KF�� �"�*m,ɼ��S��o8���VX�`{#��Hȡ���;������ץJ��?0dG%�F����YGTh�۩1LN�|^<�$���u+�e�6<�N��p�i3Q.à��4>�G�`��$k�y+���\|&�x�Y��n+�9��-|���e��=�X��	�b-Y�bs��5�*q�:��+���'�
&�!.�AAH-0Xp��rDn��>�� ���V~�i"�}w�k�c&�ל�܎�[j���7��h8�!v#����|g�[�����;/���)�L������c��ݔ��_�F��d!��p�ײ���`�}���h�\��V6�C\󙔶�W�}�e2��'�6�S�+@E���ʗc[���t+�9�v�Ѧ�MW�e�É��q�����?	�)��k��}��M���8k.���s�I���J��&�>���Ț�Y[z�|	��g�ۍ�?�&Y��Ҋ����*d���mm��w���s
� P)���Qɭ���4�ތl�P�4)��^w^�0����7����ĵ����WY@a��� ��L�9��+&CWY������:r��(�."䛠g��:�[Z}�j@�	d�A�GC��J�Ff���v���"͌��W��#�����7*U@,�v�Y*��R3�@��G*p	lM�Ģ'߻{8�}a?	��W9"-9D�r�<�7YM>W�C�G�^���Z�ŕ�zyU��v�2���Oe�N�!�Dx�dݪ�S����IT��ǜ��P�8�/|�j[�zfI7g�qDg�D����a?����ւ��K�
�;فU�������8�'�j'l�a���6d^:���g�it�]��%��'@kc�qD�,BFǶ(F�j:�a�=�bhv�㭩8:�p%�o����Uϖ��2�V�^��ao�~� ���;҄�:�h����zZҎ������˕��}����E��79�(���2���x}������'���4N���Um������"��J���8;#o�S&�	���h�E����[~r(�!l���a������ꚻ��R���\2�~"#@��qE��R�e�K;�Uj�VU�����;��Ң�#* s��d��Xt�����k�h̷�v��8��eI�[F؍M���=�jI%�gacӽU����p,2P��>�4kW_I��^)���gY����%F[�?���Ě�/m�)��^�p�9
pZ����l�v�U��׫W$<^"��VQr�O��Q�xP��ٿ*j�5��$_��r���*T������=�C?�yz������,|���+����l/�"Z��hS��R:����M;<odq��x�۝�$JgTo�kᱳgcR�8wq	�#�$(W@�����C�K�郂���9�y_�����8lM�L��6�b
�-U7����-��y�9F9~l �j�]���X� �$&:��Y�ӹ���Y�~?�t/~��~ў�]")pN<+�M�B)��:����?3���{k˾��|B�Ⱥ|��n��4˩�$�9+b�/�Br\C�yOzyS��ڽ4��ٻ������F0HN&Y�M�$CE*�Ѿ�+ږ�t'-�vo�=ҧ]σ˖O�$�-֞�{Z�#�'��7?rL�Ju���"�	(�r%��aڦ�c�\����I�K�2�� �W��8H
���:�_�M���R5mva���GY:����(쾖��G���9�9g��Lx�z��eF��b,~��Pj��/B\D�_�.�`�%�'�=P�#�}�c���	�~pb�B)��5��sH�/��8X����$�KS>KF�8@�MA���9
�q�S@
����Yo��c_�t��e*d����~�^��*\���=_\��,���(hS��M�A5�g�d����_���I�0Q
��C*���v��1P�?���~�H�(�?�Nh�[��4X�6ԆR[6oG��P<sm_����	�S8U�]e�2��d�LX��u�!�`1F���SI<ێ>�C�S_�Z~i��rS����*�@���Ѷ�Z�ԍ\g���җR�wd�#�䢪�$Q��iG����ji�}L��x�1�|V�Y�.��߫1��J�a�}����I����q Ȳ�T���K�?��~?y���w	�׼��n�����=2�&W�������QqXuqX=�V;��[�pbe���L�d��3����G�D���NAj��`Ai���8��x` ]雬6�Qkm~��	o?��#1^��;;Z72>���\q���EU�%��fL�āFn�R��P�/+� 6�����p�	,�H�B�-�y�hQ�o=���w��A�fHvM����p�����JBI{��ŉ	��y��s��e��ɢے���Kvg���e��q����٦;m��4�]-��I`Y�6���[���ܦ�%h��5�R��Fl�[�e�g�&�涂Ct~����2k�F�չ/�)>�a�qY	�哠K�?�������lY�s-��F�J�gy�vS�a��3$bX
/��4�76��rș�T��w ��t�Dd�XlxV64EB     10f      90�j_���;��l3�ގ��>�Y
�ɷ�KG9b�%LI{������pY����5!^[����p���aV>������`��i���"�����Ed���.�d4:[@>�e}���c]�Ѭ�d�o�vƋ6X�:�E]�Π�<*A�