XlxV64EB    fa00    2db0P/,߯qG��N�?.͎A��8%gNޚ9�{��<��P��aU#f�@7���[�$I�n@��.ɩP�ܡ$l؁���ԣ���*�I����,R�h��0��V��~�NƳ�p�̀<%C��4jN�v��u�C}�K����΅��Қu�%�К��(��/F g>�^I�5����#٤� -�������x@�vVݬ �W�9;f���������w�N�jQE[���>~:���d��2ރ�#C�߬��S'$�������m��o/�A���i�`$O.�g~C�L������:����_�?�v�{5X4ƛ"��I��J�\�2|65),{_�aF��9g���W�O��y��:j(�Sj��Zz4��57:�G�!~��X.PITv��񑮸�-�R��Ŵ����2�M�3���08�g�ٕ��ttx��������� ,��'r��,3�T�D�O�a2�A"HT�`��oyllVx���(Y���>(��B�6	8`�]�����4� ��v5!E�?g�Z���4��~&DpO#��/@�T�b��A �JĨ���Ơ =�h�
�P3�I��Vf�s����u)a+&�dK�ùo�t_[�m�zP�)�l�;~������hj����ė#�P�bʘ~��DLw1v��ۭ���P��G���dGm��5IL�?X;�yV�iNeM���"�r�S�%��a��I���ų�탞L��Y��pDy�ڞn^�-�]w��C�P�C�HW�����#Hn��.9ý���z�ȱ�[�����^���UB�{��H�p�N��V�@l|�,|��R�\�!����7��)��	���ƞ�p�{�5�}o�!���W&L�_<z�s¶ ���)��YW� �y��g��`��<	��Z.�+�1)��ݐ����3������<�'��qy�����5K=E��eBP�8�Ʌ30U�|�W���HRT`���O�\�8{�H�*{Y�]T-��t� ~착;4=ە���x	W8~�hk<F�����ҏ��u�ڒV��9U���0Z�
��*�1�_������ä%&�.��'�C����k �?
{.�]$�s�뙟;/_�����ZZו�)y^�?/��d�1T�[��d�ݸ���K(���}��+�5��(\���d�@	,x9LH�Zd��i-'9FF�oF�M3K��~�^����$E��$"i�tU�|/6�]��C��/����%�:���r}��ؔ�߫��C�I�(�)J
t�E�WH�W�7Jdq[ȸJ�2�D�?�ص�{��&-��j�ʥ87��ɯCܲC��g3&&v:���po��$�"^ī�$:ŮT`X�˴��ܺ'��.#���O�bDsa(�M�1+��e5S|ɷ�ʷe�lt�M��Bނpw��� ~z8J#}���������݉��Ց�O��K��^�;�C��<o�^�{��m�o���"��.U�.r2d�_Zh����br	�b������{�!�c��A�T�錤�t�PV���̤�w���諄���Ͱ��@�vR>4��Nh�� �5.Z�k��vJ�u���[<�\N�p��fOc�������`]e�Q~jvIni/��a�JH�T�GVM����c ��8��R��adڜ|G�Q�f�~��\�h����6����e:��;�޼��<�ֵ�y�	ް��"k�7hq��Љ\#�²Z�ɧF�cS�I�S�4Cإ�ZE�o�|�ޮ*-I�e+����A>��!�kei[�����L��� v��X<!� ��YצJ�f/���5�0��"����ZJ��۷�ż枾Oƪ=n"�vj�[)*+�g��"�Ϲ�6�ś� �C8퇿�a��i$��dx�(���gW��Po:;Oy��}7�����,�-���"�Ub�i�24�8�tn1��9�Ƴn�s�LN0��6c���0�<�z�3V�1Eq�ȎQ������
Y�5+�Q�p�O}^|&���,���o"V�3`�g�۹��'^�6��W�X���(�R�2J�H=�H��מ���RS� =3ĥ�(��n�[�C����A�j�mp�W)��a���tN��[����kE���������L��%X���j�-Ǿ���5&��ъ�]
�6���U�m~���T����.�K�}�-H�f�0��ީ�	8���	
��S���%d�!m�q;U�$�$���>�2�`�S���4��%X���:[
�z�y�{�*����C��>� ���}7u*9ƚ�톋�'��߂��J�i%;`���9a�(���;��@`,̈́��rg|��{������yzlFAbV8c�+2�#�A��$ϥ��&g�\��3.�LžSyP.�%]C܃䳆�06��n�c`�nFnR��zFe���<������J��S� ���:r�7��@�&��3��G�)�� ƌE�yI�)aЅ�׊�b�)��#�����$#Q�CE����a�[����a���L>���T�tZ����c����b�Vt��/ �B�J�"�;��Y�rO���se�>�."L\�F��4���}Cy�Ur��o�6���8����Ђփ��C���7�1�Z�V��^C�'�5�  O��1�.���2y�p�W��P�O�x&:���{؅U_� �p(ۣȥ��;���К�.'�W�s8 (
C�u�}'��1-��Z	��]h�&ejA�?*s,r�2A.���F���}/�Ye$s���
�I7y��:���8i!����_���ltΪ|�a΄ɚUXᥧj]��W���FeY<�v��u��Y�w��K0��A<WE�磚�T�9��s�H� Z�� ��W���9^Ve��Z�N�c�}�X��FF��`韷~�
��d��6�?5ͥ��J��?(ѻ\nJ�4X��z��#ǉ=VpC�iI�jh�5�y�^Qu�b<y�U�w��ƞ]JB�Yo%�>�)N��fp���n\0�I#B�Y�[T�Q1"���򱥯��q2c���v������.�[w��Z�X��!.��@x��æ, ��۠=	]0]���1�x����N/��%�B?�sس�I�L%fl��4�����%�ğ3�~ua,��~*�z��h��-#�}�1\�e[gV��L%ؽ[�qI�_n�C,�k'��90s�:��*E�h��>:���5�-��y�SZ��ZMN1�QD��)�.E��� ��X9x�c���������@�+#h(��b�mz$�'������8e00;ՀH���S���1�C�Q�g��o�L^o��nO�OL�4@�����?:�R6/��~�D��X��6ɡ��1���)�u��
�e���e������>�g]k�r�lS��]�A�<���"]���^����s�vZ�����ȢQ��3#'��� FO3'/N��#O�J��Sf�L�T9���d8�����	Ω�6Y��pv��1��*za(���>oU�L�FP��|0�e��v"dK1�eOl����5�7��<��t�b1е���u�3���$vBRm���&���A\�3�=�.�-���^��վ���N�x#)�̻��Y�)P��*W��R/+�N����j'+N�2��VJg�y\/�tufI(����_U�G,���6�:�#@q���v%������7R3L�T�X��;ڪY����Z�52���h�Y%�*����S�`<^A��׀�]t?hO�!���]����\,� 3���Ѝ����)�����X���wN�<�����W�:EPZBl)|�0�l&�Ԧ	�R�`�,���/��7����xv�}�@�m}tx害Vg�
I��eJFv�Zp��=�1/��\g�q�͔��xhnqZ�ICl?O�m�i�+M:��F+�;�o�*`���R�#����ϗ�#�px�4�����Ƭ-g�u^��Np?�b�k��U�#�x��QB���m���T=�|z�9��{�Z(.����� 2Z�n�+��:��i�;R�(�kp��>J3Ro\(��%r�W��Z����۾BS�c� ��C/��)���O�sΈ�K ��Β��̢j[����>�5�s���#U����J�|=�����r橄�<loٗ=�������Y秘s�>k����~~�6}�S�-"�o3��W��ŀ#�!�ݎ�ؤb�<�Leц�Y�x�F��1DZ!�=��ƫ
���-�N���#���a]#�)(��i��$"���J����?�n���� ��K�*ݫY�L��j;���I�?�=ӫΞ��.��ޣ�ˡ���X�t%�lf�-��z�!��*8�WƎ̤��(�f����T�S��4�ᝁj-�-M���Y$�������[\<�[�:��j���l�R]XB1������D���Џ߸���3��A~�\7"4�����짯ˬ�y�i�C���6W"��L���FA�տ����j݈�B�%���$�c��O:����.�%��,aPR�l��h�`��\�{��lg����n�O���>�	>�0�F�E�ЯN�^�R�ۉ�(4��\W���[ĝ�<�%�Aq\�g��B�R�{�,[�i8���уΞ'7�ط��p�nm g�H��F+�>�;A!�[��%<�{D���$�Ϲ�`�������"ێ9��䯽K��7k�D]�!� �Ѱ��]ĎҦ�
�'�.E��a��������ǡ�����U|�Q�Q��χ�*Ss�a4�m,��y"�E�i��c%I�R\��l�SLԈ��S�� ٖ���X�r=*�]Ğ@޽���8B4�"'t�]�W����o�%�n��	v��0��X�Z=�!�	�s�c�42�W�;�/$?��ܸ�>?R8��$�!�
�ȿu���Z�����A�í�t7/�9��a���@u�׶;��)Ũ�"ݗ"3R�M3�8=�(ؙ��cM����?s���� ⍴�Z����p	%��4��^��
E��З����`ٔn��Ҟ3���O� ���V�T�6�\`�K��N׌�T�;j��U;���?hw���Y�ib�KvScN3*{�4 ��^	KI� J8'(~�bS�*4bs�V��#�P�e�� c��5�oP��.?�\	���wju��[�BEL3��xJ=�<��_ѣ�+��f��Э�M�K����1鍺��t����l}�ySc|I��r�e0��6��ւ�/���P���Z�Y�	�M��7m�RK��X��"n�]%6��w&G<��2O��c�ƿ����|�jl�p^�G��+�g�W��Ʀ���t����x�6pO�P�R�խ����LJ|��ss`�J��cgi���^+���`��ded��i+$�
�u>�N�	K�����s7ވ�q��Z3%~���$p{p4�0*�!��D��i�).�)Έmu�p �ݫ=��@��I�|T*B)!#���6��n�t|�ۯ���s���KA����u�2��P�����&9� ���-?�S��sC�x\��g���z�Yb�_�o�o�Ueu��E���^=.Y�����u[閻�-��sX�T�hycȮɞ�<|n=(��Ҽ�`�����)S��G�8y�c��M�8�����	;�0�� v
t�L�oV�
u��V�t4> �vde��w��ɒh���ן�����ɴ�M9���O�*��&(1��AL�!C	�wks
�p����������mC�H�7�����Y4hJt6#,e6wBNC��H2��sHl6g�,������Y�����4>��Rʳ��v�ؤ��,F�8�='?�L%y��U��]<v��l4AU����(�{~~3�>*�ػ/�8�S�DC�@�`dx�N3\�PL_Żqvҵ����kw�Zy�c�'B��Y��X��e��f3G,��n�G�L'�ǡً�c*-��0o��׌H��Nbxx[}�'q��.-B����J!U���R�,RH&�J��[��"�U� ��˹��݉����<�3�&2\-ͽ�Dr?�{!U$q9�'��U	1^��A���g܇MHYMX/�uk��������M�C�\�`�W�R
���vj��d�;W���0{Yl�B�k�(�{�� 4�s���h
wf��j.D�������6�! �!�<j/��l��^4*.He�������P�h)$�1H㔁��;
f章d��7 y��.�f6�w���� �S��]��B����U[�!䈎NIO����fJ�/c��[�G{hnW�p\��v�y"�h��&��}�ʧ��op����:�P�!+M�/Ѡ&"�*���U@A~���H����ؓ��Y����=�^B ��1e��p�����_����r���Ɣ�Z��\�2��� �w1 �E��'*o%���5e{�Ru��&��|��n�֓�8�0�j�Z�|Ц����jrǉ�~Q�jN�q��@Ё������k��; �����x̠"��W|������+�2�m[�����⑇���S�I�BJBd�=?���dv�����AkW�eW�!~j]hIw�@X��XT;���ᦸ�sm���H������q��r�K 
���U�c��.Pj��A�&o�3t\�7![G9����8�h$	��;��RT6w�=B���(�A[Lr٧�3�4n���jp��J���w��@�HA
-^���]�������3����T�Eĳ��:���h�J�AB�(� �C��:�5�9�lr��8(R� O�+X�f��#�6Q2A�i3s�XS_o�9n� ��m"
=g�RG@��`[1�?�_)��8#�j�
� �U=��7���|E=%���_�;.�j�LѼz����_���kx�Y&�4��+����
�ya0���̮t����<_;ZEEY�����s��(����?|7CMq�>BT�*D޺ѣ����9�!3���j���J톊?����F��EZ��D�ù����%�*8��<I[�>��[(��1|����~Cۉ򻵎R:�����;�W���8�v�}��'�N¹Vw.G�<=�����QM��T1����_��0�,��i����!���k�Uc�_��B��b��w��3%q���Vj�},y��1:���$EyO�aG�mH"��doZ��&��Tj��P�2�Iv��<^�ٸ�j~o�v0-siwU+��r����Y���V�Y��d��>�!T�����6�F�=��S$�|� ��,�t RT���?[� � s��y�[�}���Ă���
����D���e��p���C��âϣ7��i]��)foH�nӲ/��b��	�be.m���H[.��Ѭ
u�.Ԝ��^�1r�p��mN�ܶ��,����.�2v��'��T�ٽCL��4�w�|����_*�%	t���Cr�������]�����Ê��ʬ�BJD��uJ�������,zQT��t_��0A���ECt��8J���e��pZ6r˩��?j�Ã�C+�lk�J����J+alTV��0��
�et�s#<�K���g��6xK�z��#9���N�d���72ż^qZ�|��'{GǪ)2ۚ�@L��l�*���P��(��U,6�(�'h���_����q̔:6�ry�	i�a:��	�D�uӧ��Y��}�o�saX�T%:�}�2}��*�E\�,M��QOb�p$Hܴq�~��s�T���W�X��v@v�[���_
�;��{���^F��,��9�:-w_���kt��3�~gwy`FFK0��Jn���M�KL�q���A��u�O,�|h�g� b:do�xEO�c �����p�{k5������ V�@i{�h�F�*�  �m��hjd_Į��Q�ﺒk�"��R^'|F\? ���=�`�B6��/(ѻ�4�ɵ�C�|���ncI�P�g��fӞ�TQ�f�>����d(�-�)D~�_�Z�����E��:�?]�3�S�)|1k�Z3�xK��J�)�P.��|av���A�H1������=u�q�m����ζ)�k�h���h����M�r&����p���I�(kY�/��36�w�ćܠu�I�~�y�@���G�U���k�<��w��3�V��u��W����\�gAi��Q��l���=�����_���{$��M�En�j~g�oOP����[�?7� L� �>q��?���b�oC3���,>3��9n3,�[Zg�r�>\�PBS�����@�&BT�\�B�c����qV���V����2
���?�>�f�Tp��m����5��DG�j����EA������+ІrjMpK��?��!s;��F*�1|�O��
:�����<@P�x�R#_����'I9�:Q���H#�/<4)'=��|.z]��|ն]2j������5���6���C��Ѩ\��k�Z�n��I
�˚��o��U�mi��9L7X����+�~���NSע1]7d����n�����q���ax���#L�����	�t�z��1�+`\�N� �{?�~�݉��{��b�3��"��,����
"��~T)z*ގ%@�^|���u��S�QF)�H������H>[dTʋT|j��kd04 ����9hr�VJ�FX�;���+9l�^�ɼ���+/��,��u�G��<�+w�5�J:0T�m�~�R���Xւ�'�wXG�.�?�0zW�Ul�2KQ��ao.T�� ٚ�|�x��H�O�I�>7���Q��ӆm�s��@nn���������ζQ���yK"����gs�� ���~�
�0���2���h������l�z���������4eʃ�n�%��L�(���?�_�3~	��Z�J���[��r�.IO����r�b�h~h�mm�w��>|N�Nj+O�*n�H.G�n��G����j��qj�� ����Пg�D��8y�=sU`Mz�I���| �~�X�	��%S��ү��b�$��;�}my�^�7�l�Z�wnv���?S��-��Xn
���x)��4�)�ܑ��%x�űZ��ᔣb�YS'�#����M���X��z�U��!Z(6�Z��k�}ߎ���#z��a6���a�ɿ�����t�w�� ��y�aC��flR�|��r�d&�4�[�'E8�q��ur)g�ؽU�ғ(�WZ�RNW���L(�󰦹=n�?��T�x�7���9�+���O�K�W�t��4�D	Rn+ͩj���m8��Z�~�m�$���r��r��N�� ���
Q�!2$�S�Ƃ�<mr_g;n��
�=��T��In�l>��:$2P���7w
��]�<5��XP�|@c���͵��ɿ)��?��=7D8�=MR1�E>�s�G�����U�8z9��ۚ�2 ��Gr�Y���2��F)˱ �y������&}�`&���z ��oQ3{��Z�)S%&��ԑ'��N�3�P��H����5.�����Sk��X�R�Ш�L��5{:���F~K�3��b'�)3D*!�;t\R��~��R	!�J�MN�F,'T�[w���l֚M*����Z�w���� 5F;��tS����*L�:#B���.�O�2T(2�rD��\�0O�Q�43ӯ��c�b�ˎ��p�-b��B�R��=O0K2��-�n�
"�j;�����觔Zƅ�>�j��LH�M5wɺU4�q
�AǞ4�B[{y��)�E-�Nl�1^����o}	����-7��(&G�Ǵm"�?�e��!vd���1��3�Oոj��º�J�D�~Yx;��E��Cv)�j��������OS��ԡ�+�;���;�pD�+���m^����j��9��ݔ�����O,՘�L^�%9k�W�cN�N��Հc�>�)H���U�`��P2h��9g��@��hƺ�5ĉ3~���a�_�t|���Il�G3�ӊ�^���wq�`��%"����h\R���G2�����wKw�v� ؂���*|$fƦT�G�ܓ�5�L�)�L�x�n}'�t��n���0�����?��Z�}��>����gcB[�+�����	�x!?9?H����~T߹D�4��[�7�E|}�"ۘK{%�G������M�t2!~���"amMV[��[h
��>VN6zs����=:���&��_ ��&_�SM���>�ʺ���sĚx!H3_�ط���L���~uL�G-�j����D�ذ2�M��4|���P�Q�ƧeO�Jm���_�@��N���55��)MǷ�-e�;%OMj��O���\\+���䁙�xR�t�d�jlo�-.�D3���A��F:��Kc2Vh��T����#znY�۱�9є�&�s�E�F���h��ޏ�t��A�����/+x|�Z7����)��p�ύP�w�'��ҭa�JlT�Dh4N]�-�����0^y0��B�x�vT�ď�s�:Lքm��s�,J��Rsa[�y��Qy��C�p"��Ь�Eʙ�yi����O���}H�XT�l�����)���:�^i�#���S-���z`<����i�����4s��{C�_��~tG���g�ڥ�|���~K�%
"�$ ]�HL�?=�ފl֒ūSJ�ƥ�z!�"�1��µ����64ನ�J��AL�镺�!�a�L�iȃa�-�4ۇ�]�PW����Io2V���٫E��~�e�s#��w�;�A�̊�A�3���[*��Jl͕�Xy�Dz���/K��]<��񧎕�,�(����l(�"��u�'mX�v��͟VJۉ>���K: D�F<zK�{����*�r����sgO+v��~�������siD��/B9	Z<��+ɏ�G��2q����u�s�D\YUp��_�K�n�5�w�"�Eϭ}����*����Iz6�~�A4q�Xd����*�Q� w� ����;I]\M��c� �lk#��"ɶ������-���!����Ӏ�R�΂
��gh
ʂq����ļ�+1��chS�s����{�����
��I�w)/'n���1ate��/A\����`����l�C���P�����C:��� +^�s��I&#�������=��>�~�\��Fm<�ԧ����P(��~X�PF�Ԋ�H͇�!x��R]
��韯f 6�bo:��2x�ޕi�T�p�����a�-I���,Z\J*'�H[�»�M4*u�9�Mg�mz��/䅌��Ua��l��d�����.��!�e��	�Df�Cߥ��2r3u)���I�W~�D��A�;�f�@���ƽ��3P4�Loݏ��<�+�@�ԡ��꒠�r���'�Xl��ݑ��*0.�e��>��ܿ�6¦HH�&V\��C#`��{��R�#�.� /{4#QV��_�k��i��"�:�:ٯr�2�uwI[�MA"L�]���6i1����g.��5�z�&9��Ï�հ1=��δ�~udk�,E`&����ƮD���g��X�󗘥XQAͯ��g}��d�ڸL�{^������I�c7���f��-|�%N]�6��i���ܗ��m�p��*����*�3ɨ�M�nmn�-v��T|XlxV64EB    3610     9f0��CI�
G����M`^�g�#���Ս6�ق��Nq<��������UI��c+�a�j�h\�D��� �����ԕ��B��:�;�����J'I��2=IHv�'ߔ�R���^&k"��С��/�A5@���lV�Y=^�A��VXJ�f�B$F�����!�{��8/lk���A)L4���E�C̷����-t"}D��'3�ov[ݢ IЌx`��0�*�_ �)2��r!�$`2l��EԞkR6��{�I�r��Wj�|Ҋ�bvkz��-鑇���Z��x+�W2��l��5�kj�XCtэg���+u��^�b������yz���z� 8rO��D�	�o6!v*a���Wث���HV��	2����]���e-Q��D��%���:ni���p�F���U'���6�/�:i�6��'Sohi��qӇ�&��v2��s"^��>���u�0�!Ԣ~��nJ��@S��ëgD" }��� N�z�,[���6N�ć�G��Xѕ�0�Ż����i���I�~ܳ(�yS:ւ���g3�'��ދ5";��?��,�N�G�H��xX7�S���p}�%0����K�&�kl���?�8��}��(�q/⨽6����_(?�0�	IҐa�0=+��=�,M�iQ��6v�����9Mo��L����7?�Rr�U�. o�xm��=�)����s�p�b�����f�i^�WInLcdf.X@���.?,d�]e�nה��3G��삕����m�؀��}��z<��ؑ��l%�>ކ6�{L�p�����;?18��g{0MR�SV�ỵ���]Wjܝ�M7 j4c�$l�����T���J}�+p�D������E�g��v�lya��-�a#�m���~%��0�h���/��Qr��e
��!.G��ɽ�]|ZLI�bR��d|N�)d����ْ�v�`{�Ts>����*�"$ѧ�Һղ�m� ���D�S�T����B�ur����,��%<FE�=��jk]?Ә���h���9��"۰��p�e
Q���+#E �I�jo;����9���"M� ���vS@�6�O�<�߀P��ގ���6��\��w]oJ���C��iO�������Q3ܚ�n5�hZb0Y�'����?'|�;��� a��|�4_ C6�k��ң:����z���zq�	��V��N���[6����}�~���U�� )Z�W�cj�%Z�൛L�K|[�����p�����?vi*<|���τ�u:;w(EX���FQ��>��G*�,~<�|hڇ\k���8T���#����P����������\O�U�$�O�!=�>0kZ	���Ke�n���$<�
=;q�r�YR�/�1({��8H��ܑ�0� �z��[ކ����WT*~�u	�#��A�oR#0�;9�M�RJ��m泌�s58u�J�XᒮmMr�SU{��oJ�4lOu�|�ȾJ>bF�ā�g�xZ���b!��߃3 	:д�������S)�,����c�H8�=�}�%@��g�`��<�F%�p�����C>�kк��D�P|��{�Xi���˙���J�A����?ts�؆lN_9|;f2ٗ�����rwD��Q��K�W��5�@�a�-i��?��F����D�6�g]7�v�	zR&jDD���о��N�����U��u�]��k �"O�T����l�|@�]|I��z��������:�`nm ���ZOڥTve3����.�q�^���m��y\o��єy�/���;��t�K�cGg��aV�x{5Ñ�����P�����(��n�B#%<�޹�{�"+/�9����38���tJ��tO��u���q櫲Z?�o�a�X�2��T�:0���)�L\{���NoaWc��hۆ��G���ʲW�Z2^�D��˼o�䤯weP �� ��q�P��I��4$To~sG�0}}�C���y&/X,�^��!�O��b��?�ܬմ	�t�%S3�*�LaY&A�[	��.�<R�bq4�z�d��<��P:\�h�"��>Td����!7�t��Me���2f��cV�\�
^��[��u��_�B >�+=�io.�%��?�4�`y�d�Eb���ԣ�����nY��T?S�jt�E�Z݋�.x�#'�a!�`i��B�����Y6�ɱ��5�^��4�7E�8S"V)����s̜�vz����t9Cot���I����]�8MaH������n�i�6ߖC�3�2|m��2ke�?��3��֕�`@������0�c��ţ��o�5&b��#�1T�+0��a�Q[��:��5���r�����-�f�1|�6\��.����Z�V~�y`��/�oc��$���hNm:b|��{|w��V
N]Ң�8�|W���~�9�% ��JP���C�1���;13� �u)�\m�΢?�z�q��x���,�!J����O�����H:brMR�