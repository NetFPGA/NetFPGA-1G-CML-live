XlxV64EB    8a79    1520�lfj��-nˠr���i�Ӛ������D�Z�)N���2�����H
�ru ��S�k�� �m���<�ֳ�4��	?�.���͉߈��۔8��Њ�<��g0��~"�T�^�]�*�a��+�c�~!��Eλ�����5��0�0�U���c��@O�6�X�/��~X��7���d�(���h����C���y^��GY�]Rz�<���<KM/.5S���O%c6	���3�/�Ε�,���@EO82�!�R�tuY�.�pK=t�f� A-J�&V��H�͍=D�$��g��虄���+��}�+�k��@Y�8�x�ۺ��O�yOV�W�$��~|@�� X���4�٣fI��܁Y���
x�E^��i�T���Z#ڭ���Ǆ�<6;��;͠��'D��e*Gd�W������[�݅�@D��n��lᣧ�O��.�3�I�۰��J���x����)R&��j �U��L'e �����w�\".�2��RE�a�*��(a_�1�Ww��>Y�?Y.����F_�����F��5��L�Χ̮�*k�7gH<6)=�+�������C��Po0��9[^�ӣ?�p64�V���6�l������b��\> uCP}����S�ʈ[�9L@�����H���3�B�Mr�}2� 'iI���kN'~�'�������*�*[�0�FR_0�`��Oo��~F,������ލ�����Ψ���U?B
�h������[��hR�`Jw2l��bTٝC�M��ƠO��ة�1����_�O�v����</j(�"�7T]ݬ��.�)��h�mu?�8;w� ��$��~�c-<��%�b�Q��m�4o���Ц�&鈠�Z���-���.P��?îI7�|?Rǰ���o�QQ��!���maL��F��������/����W\%�4��		*c;�ဳ�/r֍����3���B�w�A 悸)���l�M�lCђ�yƝ�����s*���Y'`�����.C��6����ut&�Mv;8�����i��s7���LMs�9���IW��RZ��t�[8j���o��q\D�ʇ�!%�9��߶�.��J�`����7T�1[(���zj���(,��@�ǼO4�$I�ךșRܾ�0�pfy@�����?�L�Bu5(b5z�{6T9���W���Pн�-"��?h��	K#4���ߦ��#���x�����'�&�	������@9��EJ��TS���\��RC��6����{��>��.1�B�Dx.U�P禅�_��Q%0�V�w��k[K�D��94��Ӫʪ"b�j${-Ո��m��IVmk��ET����X(iK�����::��J�JHP���l���[	Z�𒄆����b�w{��Z��
���MF�Ћ�a��wS,�&N�Q{��.e��
"0c��y�;��rHDT��F�����/$<cՠg�s_ǒ�J`t����xf��~����4&���ȚG�u�[�JM{�h�_B�r��ձq7,�T۱~]Y;_EL���[�;�a�N�b��S���࿧H&O���B�@l�8�R�5FvTUه�6'��<v9N��g��a�c)|%ޝ&!�瑇��iS7�?��\9�׭nP�mVZ]��Z�T���o3g]�/��eB�'.:E ��p��
>�A���偅r���;������-¯RHn,V`�n�P=���*�^��ń:}L�{���ر#��-U] e�,ʅ��E�g�O}��J��f3��w��(ݲ�=��}Շ��o�C!�+Q�E��'|��V�b�n�j�,��)_��視�^���s�A���Z�����w�Q@�w� 8|ZJ�v��6�y��ڒ���(�� ����9��Yoc �ܮ�w}PꐒDP��I�ؿ�"Ƥ����5^i��]Eޢ"�$=f����\1̻6s	.
����%U��;��m�����T��L�R(��+z�bÈp:�\^>� Wu;+�Ԍ­��V��\c�
T��L�-,�)h��V��f�ô��Cu�D�/��q��P�36�{�<ꇁ��Bҳ���	/��)'�:R]�U�Y-/i��OnX��qc[��?��Q��-̕��G�1}>T�:f�w!�1�SS�.0�{U,N܎�p�</v �}�EA��| �6���Ş�A���k?±�G�HBs���� +pz��p�X�2���BG���0���4w[q���֫L�ⴜT[���j�(昵1���Fyu��]Ɔ�˱ٲ�3|Uކ�����tR���u��p�H��KK��X	�U!&sZEP��"�ڹ%����"E]�M�	;�){�
��(��(�V\�ljɱ<w��&3A�-�X��I؁�9#�΄AD�خq*���g��KT�h���gU�q0O�hC���˂�+H�J ������[{��� ���7��gQ��<��v̐�V
�]�J�ףR�xÆ��s��-���!Ս\u�h˱���DYH�4�ǑL��9���J2ć{����$���֖۰E�?� �H??\�z�@�Z��(S��g����dlJ���K V���V�j�f͂���C��o�H�����<ܲ�WB�K��O,:��wY����NO�O_�T�#����MOՆ��`������?��(��@@+#�����*�~�iI9l[{vݩu�*��P��Mm�����G����Gg9�V�o�R��;ca3�z�]�J./���sOu�P���R`V|�Վ��P�^d��r ����\ڡ\@�r�X=#(�'����'��Z��m�۬�S���v ��8??��y&��0}�Xy<���B�N�MqP�ReW��յ��7��=�S��r������Ǽ�91��lP/#I�n�VW��v��ep9�鲤���gj�/?ګ6�ЂQ�dR<�g���D��Km�H�H۴��O#t��C�����}�K�[+	��`�qna��E�T�E)�m��Ehs�����ن�l_�`o֤���^����8�cfPZc-ߦ�����\�6̄o�8?)��؊nF��];8�0B�ȢR�e���Ew����#�A��7������A�I�����m".��ꥯ�Kw"��]/�}���µ9o(�>d�t�a0o�i�0�0�}�ѫSKxE�Cs�)��mD�>��܈�_����@�~�Tp(������^�6��ID�/9�QϧR���͆��������v�5$�q;V�/�3�:e9[�")
]�ZC���܋t���%�����a;M���\�w�[$��0�����Q���\����4��!�����ȘS��U�b�{��ݪ�n�kl�3�Q-���Ir��X�52S�:�a�m�&(��w�KK�N{��Ŋ|r0n�V�ВsM�
��w���=;�70�ȯ�=���%�_�('�����E��;������ǳ S�$%C�v�K�^�d����9s2�׀�^�L����S;k��g½W�	䬖O���u��p���DM�{���]R-`K���ī'������@������W�c���7AO�"5�3�{N	�i�Z�r,«z��cc"wc�Yg�����1=�/ts�vZi�$x����� H�MVm8�8ߚ��e�tG� ڛH�	��k ~���4�����7��t�v� >:���}n�Z��˻���ݣb��I�\9���阑���#�Fu�'�'����`���ۆ��*;� hn��i��.�ܶ�q�\���8��Z����������ݜe�����!��\Cf���Lv�3�!CeY��t�Th��xê��ܯЛ��O���(DǠFOK��q`qdj�:�UU����V;�a��E&�<�Bк�s��vI��I��}ʹ�9�0u��8������7#�mf������������c�s�S������U]��:	�)%�$���P�Y���QT�\?���(h���/Ѐg����=����ݒԳoǐ��mue�.y���!����C!eDy;�-�p����O�W�`�fG���&ߘ8����c�E������[�p�F?��հ{U_Xn3n>��Qs�ɴ����2]T�C[+�/�����2Vx*ﭑ!>Uo\�[��	q<]�^8�u�ӟ����Za�Od�}�ߞ��aK!�G�~��=?,	8z
+b3e1�b�o�Kde=ހy!rr�� 
�l��;ꑯb�\Sٰz!�.��#jf)W��p~��O�-��S��?��/a�J��;DB�υ�2#(t�:�[K�� ����Xz\L��D�*��,�"!R�����m��&~��g�v���=^�+}�vٙ/�'c�LAsf� @X":���:�4���-`�P������ZF8˨��>Tz�T�k�I�yԝ=lo�=������e�/s�@�|�3\,���"w�qr�e.�!N�� ��zg��'�Ll@:��o�Uj�}K6#�~�B���䇮����4�LO�K�9��|U����x�@n���˵ݦ^
�����{�qڝw�@ed��"�js��T�8Xn����5b�ܠ�����4�&�}0�C�Aԋ�oǭ/����V�y�����i ��?B$�S�z8"�љ)&i�"1��I����87���S��I=����Zצ��O�R���j���h]��[��[�{�PI�� �Y��GMu(�&PN��T��g��d��2���1CJ�8��2�MX�.��P��U���_�f�[���?!16������Ʒϵ���}�=�j8��	��G��m;��/4��sN��΀�g������ԅ����$}L q*�	�����b1�	��5;k������r��p��N�y�����m���
'�$����b��${���{s_���� �u��LJ%�����N�!GǹrG��������$���l��#Z(QwwEwGd��b��!���4��N7�;X��`���_���z�9����7��Z��*h��ҷT �s���H�!PCp����Z��ZJ�6��V���W��� .��OF���~qp��<|��2kb��-����X���y�[Y�Ӗ�UHG�KMI�^(������w�ɴ�j��
׿�}�� �R.�bz���U�Zzq�:|���y����*>�B0�k��ť7�KZ�>�ρ�@��/��1�/Y��Ǻ��N�Ϳ�|�,
��-�!��9�d4�X΋{[�X�֨�h�횔���������|�KT�E�4�|����K��u��M
v�!y����uU_��b���`�80xa*l��g��%���dn� /y�'�DW�Gr��C�
/=���P�ȉ�