XlxV64EB    8214    1470��N"�KZ+X��R��$}��SE-�
�#�l$�S��f��%�A�޿l��Żv���G([/3~4?3���\���x���Sp#�X��[�&ǒRK�~d��|g��tW�N`y[+Wh�w�_Ou�����`�.���*�^ɸ����^'�}��V�U?�T�"�"�P��|�N���ʧ�����b�wK�P��r�杙z}���jʪ��Ӏ��7#�6�ؕN{��_�O>���.u),�V����ό	!�>ԉ�[��j��=>A�0{xF,��g���H<��⴬i�l^w
z��.��8FD%?�NVW(�7O8=T����c-@[b~�q1��NV/�7>���j���#���4ps�`Gݤ̵�	�6�[q��~5��7�@0F��B�l��x/Q�(@��Y�yP/;��?�E59�7�L�#m��_��X���Y����D�pm��SB�h���1z,�V�MM��Y�U �ы)�v�E��6SIq˺��R���a�ʞ��*נ�ni�9F��W+�mGo�l?���_� �N������� ]��r���V�@�[l�Z�|\��8	����C�s�,����w��btw}|���:�'<K[V������o����'6�8[�b�L0� ��М^$�ߓ�A����ա�����AR�<
��LK��j�d݌��A"<ŧY��}O�Sn�kI�&7��Չڡ����@_t�joӰo���L���/��6�*}�؝h���/�q��B��iж
�#���������i���^��jW`���A
~�S��K�/k�`W4��y��!�� �̨������oeBUP�U��d�
�.`�n8�mq�7�(Pb�l�Ţφ��j�xz���#��b&���W�y+��my�v%
;h��ИlƷ�x�C�uB�I��Z��e�c�/�nc(���|��}��4��r�"�4�,�C�U���4���Z�|i�P ��Mm�uye_<�ƋM��f�<QH!��H����P�Z��]_�����񐏤~�j�(���v�����{�<U��<E�s�u��4]����C���M�<��ғ[:;�<e�ξ�͘h�jF.�h��}�T]�e:�G���-w��r�B��"|�#��������,���7������;��܏��A�Z������0��|���!��X��L��+K�����8-����f'��s61�,N0f7�4��ORF�~��S���ۀ��[cշ�au�
��O���.�}dFh��0c�n�X����:�&�)	Gc�̎��Z�=�W~'������V�V*�M<C�O�Lu����ʌ�+tPۖQ���/>s�.��>�E�T�x&NG]�&��ɫ�iA�'��7j*�����
x��`�߬���JH�����lA��E��>���A`� a]��"Ќ7~�g[H;��J���]F�r?��?�%"��ٰJ!��/����r�`+ŴUt�g8oU��K�7�IN���k�ޡu<r��o��$�`}F�IY���䠤2����x�%��ۅ�n)E��FJD���_Z���Q$��49��Hz;��c a�$�۶�D"��(�A������*/��gUoG�#G�yu��r�ޗZ�j`�O�5#�N�������	d�QL�[����3YƉAΊ�K�@%a��o(�kY�'-/;���l�!0�A�����cW�h��g�)w�@OZ`��Zߘ��w��V���(c'j4�̣
���n:M7 �ؕ]ɗ�&;6Z`|�6���}�@���	�4�����q	$���VF����?� ���l�5O���T�� :�g5��A=ĺ,�*,���������KR/�٩ 
�׋{������bx�^BJnes�`�C�!��0�0�u�W[�˨kE��mH���%@�/,��$�`!�C��"B"\M10N��1�ƪ'N��n��@�;�v��N,�;s�CG��KB(y�+���p�TP�<@m�;���-�1jZ_�q��!������E9��phҶ���|�����w���2Sii<��%P8ұr���,8�RA6�p�����s�a�܎$�/ed�g�{�wY�XR�,�r���X�!�<�Խ�,^��|G�ьρ:��D8��s�,��iC]�3h^E��R>�ĭ��Hj`1Fc�A�5l��$N�v~�^��`o4����~ʬ��Q�~8���+���<P�yCc	6�T�jW�@Pi�}��JH�' �I�.�Θ��A��̖e@d�%rI
��硧�h[Z؋J��@$�$av�>"��?`�_-�Q�=F�����O��/����~�u�M��|��̜�<,V�;���7�2��!r�q���e01i@���Ң��g�#�u����8g��_X���R֮���n��͏<	�
�Uۍ� ��5�E��<�~��NJ��P$�28��|毜u��0\iD(�'5t���Nm]!f
)�XUX3�	\�v}?�7ǜ���̮�v�,��o�1\@��I7E��s�t:ʂ��)���4Y���H��0�m�vy��=���IbUɏzضH�jD*��8���©2�Tq����/2��QC��$�Nt��QB�=g&�f���H�~%�t��(OQ}Tf+#ܠeNZ��)����v�)��kv��=0��1�QڮA��ʨ&���L쇄�Nz %J���jL���XBj��1�����`2(�Ӏ)��[��3)�#�\��.��Xz���ƫV[��c�J��
�o�$�6!���%9��i\��`#��MA�}��$��<lK���Hh޻.?%�p�o�~�e�iSx�N���.�Z�6���4�MW0�Sj��>���|![>�K�L��O����q��߬��4X����2����̂��Dlw݉�@�m��X��u)@��ǳ��	
ٛ����Clv�J�IY[������	�����[���Vt\���5G\4���]w�]WRyXR	���|}Lu�W��i�MŪ�_o��9n��\o�;ez�z�D���Wz8��ߵf�hM�p�~�8�5Y��L�8�����C����ɾ�i7	�}s���T�i�z��\�oW]��^m"�o��%�$��{_���������,�F��_V�!!C�`�����g6C���`0<`Cd�w:A'��|i?M�"���>�E��S���'��
�iV	8?A)N��=�����+�G�b�<U���y�����!�bƉ��
���>��B}��2(�I~1i�8�����Z( eBYA$U[�b�>x�:X����� ����g�f����f/ql�������][��Upgkҁj���D�2�Y2��x����Y�o��ˌ������]6�%���>�-�9�D��Ӈ���"ΈL��6�g� ����D�Ƒ����	u`��Iy�` Bx�A���Mp����+�gx�x)A1���F/>	���Qɇ/�ө��'մQz�q3�nY�C���)�:G�h�E��*W���-;�?.o�u��u8��-�ޗ��6�����.���D���
�a~�x�ڥQ�(�+��C�{,���(`�Y&�u�k��d�»0��J�k�/�z�T�f[����[~�� ک9��*)P���U����g�P�w�z�Ա�Ȫ��'q�M�>���w��,�����b׾�t2R��<���F�y�r?���ց � �兄��'ʴ}���'��B��0&��Ԟ!�Ҩ ;f���j:���N�H.@.X|���{�);w~�l�	�E�h�Cq�r��K$\$.����ŉ����c+ �E�rc��s��[��I�)�k��pC��%�ɽ���#���Tzv�Wnq�>����.]>� ~;pWL�f1��u��LS�c���(�9��W�����=I-kNx	ސe[�ƚ6F?���aj[vh#S��0x�a:���/S���̘�j*�w

�\���0��iFٜ��������[���x�N	�[�``�\���f$�"���7ຈ1@S4�����J�k��+S!�s��}��"5�����bu��=�+cLyP�d���\:
������?K��й _b�փҨ.��f� x]�.�Vid'k�.XLG;/M =�t��Yዢ���ͷ�B!��
��o'D/!;X&u��Huj��Bo��n���j�OL� ��ޯ�����o��I�C���_@l}J�`��z�J�IW�3r��}3v��;�%����wP���b���eh�*�h��9^~t��7��%��>�wT��ZF��[C΢w�^Zz����ׇ��|C~Q�@�FՄC�9����۱)#4��FI��}"Ou�a�~[�S'��$QO�6�f��meuPaT��0ݒ�,ӝ��O#�~R͔�>鈜�xXs`c=���.'���]��x]�sW�6j����-vZ�o�gcQ@K-~�p�u[���F6�9��%��u����s$��`χo���W䫠�W-`+`զrt��ԫ�H/��@���8����?&{�S�L��_�m�r�
�Gj%�,��BWBr~y~������)8�՞�U�Y~�� Ϲ:C@�gT.qx�W��w�M)쮳�	�0?��SG���Qz��{R9$AY����!�"�W5*��jL��h�P�tY`P�����'�f���iLF��p42���Ku��S����8�q1�z��*W��;���'�K"�s`���b�����|�m��F�nR�w�lRN5������	އ�L-j/T$�&<���1uW�]Ok�@�����I��'�Cr�Ϯ� �������V��`Ke����P6��� ,�+� *��Q�<��$�T�d�qr0�Fy���{]a8�8�cs\#,�('��GBZ�2�z�����D�KXM���%2=w}[�s�p���_�u�c���gi�2��pD�6v��V��)��[�2oK��EOA�U;�>_���u�	XgX�pü⨚X����} ��x���� QM�0�|)�[�.�؋*j�����=��׳?y�JYv�#I�X�#�����h�}�-��ƅ�ݏCN�P�����{���;�ϓ�j��)R����1��������V�ku�=�f�V�*�OZ���M��E�N�Q`�ܸ���$si�g��8�k���1_�=�|2��