XlxV64EB    56e2    13e0B�S�%��2g=������C!�S� �*���0����Z� �Ou$9�i�k��9��Z��m��C�$z_���rT��L|��~���~��h�~�M^��
c[X�K��f��JiFڌ�Z��U���G�s����0���29c=���������c�$�+���o�%�A�3��6�4�Zb��}�R���W�;��E���s��������oɻt��&�׃^��qӢ��P���x�${��C+���U�B���~Z_{K
�>W}��Qw�c^�ַ`�+�V�[�1=$r!��g�7��O��r��m}�c�>�1
�%-^����i%�#Ҹ6��D���g���boVB��(��(�YZ�&�A�����Q�ʐ>�t:6E	�ڎL��'��B̍�T%cWnw��Sw%!������n��[���ۜx�iV�ᡔ�W�(E'3�qފ��e���?��R�T�5�vT�0���j�7�ްGӈW�ծ�F���'�V͙R(zxFG.<��w2Y{��;���,�$6WjOQk���?�.Ԩc�m�yzI�*;U%>�Pܚ�,v��oG^��ex�ptϢ.^y�p{�3��*;I"�p^��#�{��o�#�ߛ��>X�\�\Z/��K��4`�����¤r�m��=��F�E�xKx�0���w��=�}�-�ss���i)��]��;߱|��0���K�n�
$���F�� `>d�G�Q;&� �O<~���^E [�yҥ��^z�[��[�.�Hd�Z5��x/�q�7A����6��nuA%���ܳ���Eb�ɭ9����vͽ�H�}�8��y����h7�q��s��c��͝Xs�E��<:.�i��[����y���f'w($$5z?C�vr��i������>LU��Î`��g�9fL����9 Ү,**Z��V7^$����{��ox)S%�LZk��w=U��	$@-R���bC�5��J�ݰ!_��hEZ��{ҥ~�TtZ�F�V=�Pa�����b��, ͗B�ς��*\�&�K]Ֆt3�P��+}'c���c#I�^e�\/1�N�2?��u�o5��sF�j̰)�&법P,�kĜ|�*�Nsj"�ŧ��������gl_t	�V�wL�5�9�H��h=M`)���u��Z���	��^���Qcb��t����L#>Ey� �w�m��,�|��S��nb5s�Y�'�rMaYK*�hS�t���:���(�%ȍґ¡t�
�Z\&�K�s�a��|�;jޠ|��s��k_Ɵ��s0�Bk�#������
oJ�M�{\�t�wP �cT���30�nY���
�(ߦ��U���/�]��$`��v�%���E^Y|1v�f�\��a��ZE�����l���Ky��~ɱ
��>��XX61@;�+�ۿLُ��Y��4�P'�l�m�iҝM���Ǝ.Z,h��3��2HT3+��-�c8�c?������9�),�i�M2���s�>ߝ��W�կ��I���w�T�j�8��O1��l��4�Т�#��y�|�u�����nz��=�8:�]O�!v�1��*�X�<�Jӻ��F��1s�mԖ��jN��|4v�������6sQ-�`�w��/���N7��2 �6�0�;�.����8�G9�A��c�~�trG�"���-�n��)�<�M��)p�k�o����{ByZ V�z:	�Իl>J~ۋ*�ڵJn�)���7<�#�߽B>p�k�9cջ�?��0Q�X?v��q����>UR(W�/�]���O��8".?_��C�n���]�2�:�t&�m���>P)�\�.*��]�Nm�����إ�[�Cs���`l��(��ۭ�8�9�����x����L��#��\z�U@��P8��z�������Y�i�Ϸp۶�� �K9���k��FDo�`�]�|

�8��$g�n )�nY~�!8�~���Ͳ$F��@�2�?`6�	������X����S=~BH�.�Fv:����&��@qq�m ̞��>D�>���#~�_�YpA]�-D�� S��J�{�̓�͍�>6�*��v8�����:���Xc��PSY㴕o�ش&�����\�J����#.� ��,2i��Ι�|s��������H�H0z�,�Vdt�" �}�R�+�>���Oi�)��}��Oa��-(��X���x�Aw����x	�+L���`�JK[��jnici[1lЋ%������!~�+�Rp��u47�y��}H�M��g��r.H�����֡ _Z�BG��f�����1�.�tk���?g3?H�v�f��ߊI�6LC�IU�Z�ª������C��~3��$�� �^���D-~oh�[F/s�!���A�	yU$��^F��(��8o������z!���)ʢbF})O� ������A�_���e4�Z���HD��Q?G��f��\�RG����C�C�`�:�ZYX�����f���cM��������������;�(jC�N
_�������@b)WӼ�]�NĲ:�q�B�7dk<�7�졞�a��\�3O]�1a�����XQеŽ��g	�J�mZ�l
=u�C4�L?��q�����'Rz�Xk�/6�;)��X�t�'_3'���s�}�U�_����8����$�6�U���"��U�nݪmۇ���	��(����l�ƾ�c:s.מ��{iN��]�g���/x���~�]���#��br���1��=O_O��2�d[募�]i��1��:B�`�|�/��YV~����\�USu�ճ�91h1zo<^��R� JhyZ���2��B�Tm�3e�n���u�-,���Ry��L�)��gL��7d29�����يy_�����ɴ̼��B9`6=R�쎅������t(][T������2�Ѕ�q���<�[ig`\�;^N�yw� ��F�x{uf�>_j��#���5���c���~J�+�B�\J_8��*�ԙ=�;O܉��t�P&&*;`1��ko��=���D#��z��k[�ݯ kh��ָӌ�CO��>�e�P$�z�<��H��]bV�(�D�rV�7r��؞���éD�
��b�ӄ�����Gp6<j�e'�G���ZH9bS�z�١!�(D�8J�a�f�
3}�>�	&�N:��3�~
�kt���[[� �ѻ����km��E,F���wK����B�Qd��7C�f�VG�yW0J�7�H�����/���C�6�+kX�#4H�u��������؝;��l�:��L&��c��-���0[i��+Y.F�o]{mФ��r�vPXF3ņ���&�d-+�}RS%bWOJ�	\�[3�ccw:x(O
��B�����(KE7��QVÌ`� O��|A��"��5Y���h�ėp��pO�������ƪX�}������[X2�s�v���;�>DF���
��T%j�e�*���ԙj�~<����g�̱�1��~ ݰ] p}?lkV���@�����մ����s	*����~�Y픥��?6�5F`�s��x�����9-�3BXm>�4�E�w�c�"����8�H��F��=</â8Iל��{���8#9#�ff�(S���̚?h���u����\اȃ��v���u	�H���+Q��t�N�
��7�R��G B!��li�1.E$$2�x�!t�fv�w&GAAk��Y���,�>=�f���Z��φ=�\�������b�[39��dV8��7����H�}2]�Iø�w��E�x+�h�!�5��IF�[[R�n.M)����aǱ�_)u��c⠱G$����<[��z6�iF�Iy��QL����T�	���z�G*<�&Fw��T��9Ēi�`XQ����X�&M��YL4Mr�"�e�@A�?�s>��KB;5�g☃�y/�t�q6�lG�"ڙL)ݓ�d���������e�D�Ј�i�]�Fa1Ȕko��_�.$��C>5��ô����
U�lj0�\�̙E)�̋欅C>��r�*�uR.i��i��������9IDo�!
�&�E�0RL�$h�V	i��v*dSTʍ�����[�1�ҵ�ȃ���{4�o�o%�����u���P5]AR	�0\-�;�[C��������_�6M-T�Ib�X�Lc�W�ۄ��yp�&g�pt��e��<����D�xȲ�lˉ��a�V��Js�.X;J��@K�5K���
�P힠��F*:8:%����x�#����R��58{�A)��p��)�����nB���vw�]��NT<i�( �V�4Ȓ�Qf��g�E@t_�cr>�Ӓ��5	ՅS]ګ�y��!�0����	\iM�'|��u'�$��c]։��~k:�D.�����)�1Z��J3+�?QUj�a���.������C+��)��F�X�O7��{��MFT�p�I�RYo��b9?-�{��]h�w(��`�Zƅ�ho���̱�� ̑�M4���[�o (�N��KE��>Q�%v���D�Ͼ������y�^�v�2����Ѧ�>�i��V��fF�`3!�����8��`��mfe�<�29����Z�[��A�&kmKxݧZ��Aӧ�����tP)�c�����\S���q+k�L^&6��o)���N�����q�f�@���́�s�Ђ�ND���ǎ9J�oP�7����qco�}������{����ڶ�v>��=��f.��g���\� �8
�9#:�v7T��,RMb`V��X�\��n�� ��4c'K�G)х�A|9�/���B��� ��Z�j�LF�I����ڻ����bl��g�G5�*��G�k��SaR��%�I���Ep;g=U*�v/W��E=��|>k�|������wV���]�� ��"5�w<?8@����k�A�[�F����Բ�L��&xF��[X"��2�zN���5��:a��3H�*���g�h.�/^"�(,��/��n�-�hV'|e4N����j���F�͌��Gd�g3��\��