XlxV64EB    4c64    1480��~�=̹�8-���7���o���[�끒���'��-�Q�����g���'��Gр��7����I]�4Z9#|r�Ⲯ��h�/��M�H}tK�.�G���*�׿#1\^�՛�(�8����û8[Eq�/E�F�(��:�]RId��s�~.���n�k�3z�&�E>��Im��8��	��֐���7u&��Z�~�^�����o���KYГ�&�ЁO�UzDC��>��3��>W���37c�D>�^03.J&�Gp՘eG0�'ܜ�a�[����c`�9Ȍ+�I$�(z%����qT��d�Y��!�1��MO�c�,��7����w����-7����p�R2V=mJW�s�x{����o~�o_�xB�4�=5�#J��U���F��DdZ�ڎdv-������O�W>"(/)�!Q�"�w�-��G�PJ�8%��ن���l�S��=e����(�f74�v�M�č�7S��O`���õn-_́/ Gn:��,?������غq�H���Q��֋���ju���1[$ڳ�҄�)/�?��>5�V�����c6�'�`y���-="��I���is���W��;Q[�?���f'm_�l��b3�)�D?"<�V�ڙ�eT����BSx/Q��i���]x9=J�(+O�������F�����
3Ae1��I�־:Ҫ`ʆT~W(��U���p�"��D����O�g5E��4Ѧ���_"M�vz�D����2ׁ'����Ԕ�(��I���J!�Zb���'.4z��rhN��SZ!�),�v�!O��~�f��3���E�wE,,��2��ڑn�N���3-�;!�ޮ�F��b7Bg�pQ���*��`���r^�����8P_�/��8o�λo`S�n҃�'���עP�y�"�,��M�W��it�����ڠE�6�Jb�^3�ޑ`DK��Y�����"��Ԃ��(0�"D�r�p����c�e�8i9���P�l��K�'�[����˃q,39��kJ����ʎ�8�r?H���>S��,��;�d��}tN's�o��_�tB^���2����M4Uؙ��\H��+�-d���c���E 	��Sc��9��.Q�O)��ļ2�~���z�c��~�U���Q��0nt�
����r����UR��U�ꯓ�!u�qam�������4.)q?�c`/�t
�?�!'Q��=/�S�9!F�#(ڔx��G[o���8��L�V�����G�h�]��f�((��ͺˁ�ʹ���I:\ޛ��*��uސ�O
TA�[ۅY��](�Y�>Y۽�x��x�f
3(N͜�2�|%�{s���B��%u1p�J:���ޟI�ί���=�]82Tv���3q�S�ƚ�,��I��z��|���9N��zg*ȼ�U��lN쏰� hHe����Ofy�:��+��f�����7��Q\�?_��"���<�:�}��*�L�A,8-H����n��S�� �ќm�"[�ԩ�}�K�B�s��{\��q�� �R��:3N�ƞ	�<�����e!�#����}S���-��O�;qc�_"T��^+$c�J6��Y"��:T����s�ܜ�5OS'����C�̳�	��Bn�H�64#�T@�z�R�����~&�*C�ϼX�����Fkl㞱�Ps_�?���``iөSYa�x����:���7"�Mm����]���%��tEw�ӄ��l�u�W�ʕYAl,�Nb�^�$<)�}��%t���VD1ie+ƿL��]�{eUC~�!�Ch��b��7�J+�F T�އvv3�7?]V�=�3y�~�`���4$��Y	;�F�uj��C�z��cK3Il]����䚘s@xq��5 ��uˑ�s�N�fS����n�h�2y�x�V�b��.!i���}2?Ӿ/џ�j�1�Bija.���&L�iȒ7����2|'�9U�-zuj�$L	&2�*�[�o��3$Ά���cg������6��^
�u�G%7�k7�(��.��E����nT��B�D�OC3�s4zl��tiG��yFtI���T��L�i~#4����|/�d�������v�Z�z�S��v�l���R��~®�]�����:���\��b�d�=�y��T��h4���	�����Yꝯ�nc��ml��z�^a]�"t��KP���G��2*��o$hvζ�G�L��Ձt�F@ UӇ���5+D������=L~��uu3��ah�s���O��v��>�cuW�z���������Q��n�J�3*j/���o�[�A.|JP�vEQ�@暛��k��L1H�:73(��[�}�Sϧc����J����h�&�چ��7=HX��jj�q���Ґ�9�k)~r�H�s��oQ�U�M
"�QE����@W��Dn:�I�J$?积oه�K�|X
��R.��25��� ��S�.x�8N�w-�<����Ѫ!��x�36�lP���������+ <p;{�@�.-�����ZV? � �I�dW$kbׂs��+`��[�h(����h5L-���Kq�8M�tI���4Dٛ��3ZY�ޚ?M�0�#�W٪���E���D�E�u~�W���8������>�r�1J��������K �-�6�{^M�~�2��/�~��]e��Ӫ��S�$ԫK��w���Ŧ[�n��� ���.�\0�&yȂ;�����չ#Pv�ʇT��7B~{�mǁ#sy�#ݢ}�G��$Ӑ�����"����X���͟M�M7�my��|�D���B��L!Li���5�)�w�=F�8�#w�}��o���\��j�hI���kQ9�Z%U��qd�wP*4�d�c^�[����X
��%g���۷^�
�NqZ�v�%�aI_�Q�D��$�S60@�[�mժ=�cV����[�����p ��Ȯ����\>����]Z���aɺ<�ڔ�d);�*^�����o�Z�eӅɸ`]�@�Q_$W^�>L攘�t��z��;ᗽ��}���?�n{�3��-g�&���PW6��:��]�2 �{��j��U��� 
U�&l��h^`{�F6��T�n������$ZT��k�5�CB��le3���t�d0^Iӳ�@�X����8�����9�%m��~����1�Z��o�Q�Y�rNՌ3�p��o��.c�+�~�h?���?d�M�
>�`֐g�4���J�[KηmR/�\�Ԧn;�N&
y���j��:N^�~�k��������$�#[�%��ܝ�L/?�֞�;2졛j����)��{S}1�.��N2Bz�l#ގK�3��'��A�
6y/[+�Z(�����5�:���O����5`<h�&XB�Nr��DY�Uv��l��`�ƫ�ڲ��ޤ��<���*�G��Ebh�]��^��ajO���RB�Ȍ!�������ϟY���TF_bp�O�	b�ʼ�{���%yPX������|h��[�Ҭ��z7b��jyC���ב��ޗ{2`���3�]Tk7T�8�_���)�Z��5�E��u�Ý�=���n�����]�����=}ɑ������y���(#�A�P�a��Р� �'���*���Uul����-9�Ys�:~_��bE�������+1}ݩ�m�4d�f���`��Nއ-�.	��*!�P��9'��|����-�{1����,Œ@f�����_ůS����O�K�.����
�c���>�SL�w�����̙���>XtO�����p�R����x+�8	kB#���YpCɬ�#���R�qU��#1̂�yfƎ.sW�1�7\𭰒��}.���w��QuM���P���}��k4=�D�:�{�+�簬��Dc]�h�f�vCx?(�!��r�8��}2@*CK��x�Y�[�t�S���v�紦h�k�v�"
%�aY�Va��tTOI2��¸�u�;�<ω%�.uu@�5����";8ލ�:�I��Q�,��[�7$�xj*�����5�FF��:xT��PG���j���Z����)>o�*����v�ij"qL;5�rx��!p�Y��ፊ�돒$�J�>��;?�S���0���s�ڵt=/�i`о�F޽�4���p$Ӆ�~�_�9s�\)F���e��*����5n~!Ȭ*��OY�%1e<@ ���N[���K�zlH"ь�ͻ�h1D���<9z��k�UW�f;��4�7�C`�F��2q }|�hϘ�<�8U���V���?c"eM�!	t�6�]j�]��ʋ�gt���~S�P�t	�arZ}q�yQ:8f�F*]��J�k9��� ���c�kS;�涅
����I���R*���z�Ü-�m��Ĕ1�l��鑍� CBg����g���b�9w�=k�}],�x-;|��_�|~ �X����@����u�M�;|8Y�z���Ms-j�y�Q
���ծ|�Ȉ���e�B�K��t��Z�iuH�7q*��c�i��Ծp�2_kp�<���<c�gk�n=t�x��e؝���O���Xk������s�Ʀ�̞�6zȁ~�	8W\
Z�j�ڋ�&�E{!��J6j.��)iK��+19s��I����$
e뮢v���Ш����O��p���~��?�-���D�x��M�����E�}Wn{�n�;3>��+���b��%+������Ȥ��O�ĺ���M7���:�PL���+<9�ļ�����N��+-m�}Ǒ�V�1�8��,f!�!a��2j{ �����a�.��k�Ȣ#´��y6��}��PM���CAA-�<L� /����vs�Ax�r(��q�h��
q���Q���	������&v�j�k�*,k�� �]l�Ez�����GO�c���A��*����>�+�R�!�%�	~���}�h���3F�������&��3v����>�T6���Z@
���.sF�����Tm�]<��x��.������J����|��"�r���)برf�$T�/e���ZxC���)	y���%x�t!�h?�D#-�l�� >wuql\�m�`�zW�j:\�,��e7������v�bG�	�����J��Um�K��7Ņs]��]�d�5jvw��Z m����