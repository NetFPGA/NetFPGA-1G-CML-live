XlxV64EB    24b5     c60UJ�?_��X�Գg&J<k{�k���;��+e�p���6'5e1��)�!�7���L�7@��W�}�����-9"�=y�뻬翭���B95)G���+���݉�է+���jη�~uo�ny�2|��:���#�ĳ��;o����Õҳ�ز�P��|+Rh�0��x���Uj�?+����e�p�}M���
^N������y&�ox_C�Ͽ`�	+�|g�\"2�#�6���ʂ�Z�4D��4��H+�i�=d5�.����3���!��M8S�q�$G�=�*����@���@�'��?y�3菱���r}�s��pˋz�hߕ�$�XoM3:�k�7�z�}PD�P�2�qAbJѶ��ɡs�[#�P��`��Y�8�w)>O{�#5p����E��+�|��q7��8��F?$�9���_U�oѹ;
�~�{M�i�����E�n��%�@���xC�?e+v
�i�
�2��*˿TQ��w�L#l�R�C�j2��R7�\z!ž�dg�����20���_�˧�X��S��b��[ʀR@�ǆ��k�Ǆ�p�c"ޱ��_��d����6 �F�O#����瑋�Ci�5%�t�;&�8����ꏯ�av��N��ĉ$�l�����+�l8��6��$i���?�PhM�̶����<웶F��U�A��G�h�ʕ2�E��I�Eu�w���\�in�R�6���.�~:>�RE��_�3��W�8�<�is�Pm��w��5o]��T�(�9�@��n�s���� �ѩS��\R ���'�O�#�H`;Fk�Z6�uU�~r+^��H�K�?��P�l�G�������]��G�����Ga3�s���PZ����� C���l�
aU{elK�s���V�>��&��dS��ᤓ>�,-�u���(Y���dś�������7�����H}��(�g�a�~�g��v슭(T��z��驱����h/A�*8g��=�0c��� q�'��2)�~�J�ib)�b�7(D~���i2�x	/\��W*��`E����p8�K��!F[�Sc�9ף\f��꼿�4�O	<JN99WZ5��@��*uuI8*��y޼��37e]{�I��Ƃ�_��žS򮋲���=7��y�Ҷ5M��J��������h���#��S8{�("ޯ��"C6J��̮��/3��ͣ�SL���:K�v�1��R�ǚ��ks����H��u����	l���)&�x驓�s��+�Յ����H�*Q�¢��
Y\rN��g`O[(���06z�ɽ*��3Y�Uj��T��~	���7:vӏC�2���a,n��I���5���h*Rp�3�g@1�x<�l��U7 ��q���&� &a��׳H��]��*�ql�xO�-��"�	��83mg����\�~��$�o��T�}�y.�gO��JTO������Ui� Cb���w��s���< ��a��Q�[��ޖ	�F�DM�$P��p߿�xK�O^�M��V��ܟÒL�y���sӅ�nF��V͵r/�y����>��J���iM�'x��C8!𞛾�a�#p�]�����qO�*�p�t	��w����ӹ!�;�9�������3y@�d*\=Qp�J�;�� =�Z�4��IԠ����C�"/�d~�<�+ߡ���:,�(Hg��d�"T�zp�ڽ%�-��ɠ�2B����58�-��! z���[B�R�1��{�|�I+��L���y�S�eWk�P�x�"�зݎF	z�.+.bM�<$��AA���~�����R�
�X}�%����'�K��c�����|�ff\þ���3O� �b��f�$:����_��������f�N,�xG���zjrxȓ�$�o}��`��?_�/6��vRF��]WH9*^�E�d��4&*�N��~���R6��J�1�)N�HѠ�3�N����)*H��;%�:���&f`MM��*Z�� e@FOӺ8�F��iU$F*�C�1_�$�4Jp>�W�]z �%Ҥ���GNc)K�l�UX���זw��5��]8i.U���)�&�����!�=�iP�g������h,�e:� h�������ԯ���h�9GEI�_�3�պ?l.�RbAȬH�*w�|�G"H^`?PP�`�X�H��峱l�?U�̞ἁ,����p�7��V,�hkl�F�>�� Cv��I?�o�j��8���	i��2�"������>�A�M�W<5�L��W_$�W�e5j�����D��]�e_�	]H����S�)���B%�C��|%V~<tL��m-t3��y��1�L��ȸt���l#[���(_��3�X�Q��!��Z�a�6��M��-A���+I��Gi�/����V��9�PŎ\&K�"�P�J�:�w_8~�~��!1�
���;:]�,^�Eh
�7R��7�	�D@�u�=���xvATyX	{�xm�^�<}�.���V$Ǉt��}X�+d�j4$��ԮU��b�f�0���;��{���T{W)��LYm���9�īKQ�60�=s-��HuV�_�9R��lY�6�tB�M�Q�+�O��Jdhi*JNOp��%��W��.9�jYND��$�i����-��*������K��'G]%�V]?��wE1l뫔�\�V�fhG�Og�[���А�]��u�'I)Ly­uЂ_��_�D,���sn��y$�ǯ�	 ��h}��a��	����/d�\ů���Rb�mn��� �����%~�Ƙ�ܳ���8��b˧ ¹0���L��WC}�~(���G<���[䢄�y����R��|k���SZ_Ƥ�-o�T̗o>S�'X�b{��	��S����w� �ꃛ���?إ$)���H��� �]�s�2r�����Y>�����#�ҡ/��~z�%o�U;@�a_2�&�r|�����5�\�"�%$罔�y�!�|��7�x��2E}�O���k9�~z��[��x/��[����Ř�P"�����N)�,���4�xR�tk�j�MJ��W�k� ż�9�ׄ-
l�^� Y	zo����+°�ځ* �v:˥r(��E����u�$��^�57������r����.8r�.���k<