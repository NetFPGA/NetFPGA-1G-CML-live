XlxV64EB    fa00    2d80u�ͅ`Lk!WWW%q��+z����P�[V{�d���Y����E��(�&�}5��Dz6l+c�->�J$�`'�T9����Vn�Ѫ9�^�UW餲�q�Ygg�	G�EB���6ճ/�!�+s�m$��Ҿ�S�Mr��>��4�v�@�o;��ӵ_��x)����K{$�Dޔ'~Ñ��z�E�#�o��ǟ�0E�_�E�� FN2L�x}��_uF7��Q�e��ĺeKw�ν�l�@�hp�z���Lc�&i���^�����wph�}�kt�| i�e�� ���t�gJ}\�:�1k����79'5YMRw�x����w�%�?�Nͨ�j���ӆP���?.�{�h��P�\dG�H�ZW&t��G��+�5�M�Y>���x��5ɡ~l�����F�+<�Ӳ�v ���"s�&Ua/���pv�-d>5[d�W�7G�t�����s��Q'7�%�~��~�W�X�̌��3��K�)��&މ�.�"~Z��V=TARl�]�퓳�{߻�j�R��X	E��0��ko�q��2�af�/	��Z��N
�*[B�zvP� �0:�txOa�>Ԍf�M]>���
�e�x�]�?ZcS�������:��pX�W�LF�0�b`k�d�M%���~7
�9���l۶j�Aƀ�{��{��l�98���=k����h=L��DiW�S#�,*��F���S(�:���T	d-/�7	W���E�eZ=���o��Sl�a|R�	�D�#�`ͺw]�0���q��uj�/r2�	x�k%�1�O=�,�Imv)��[J�k��+q�j���űP��� �f��2#��g��*���U���̈́g���Q}`�ZѼ���a�鷕}�pG^x��:w^��&�o	I�U�!Jl:N�R:߻�ۭޘ��tX�r�fDA�š>���O[������6�f��jlC�ۦ�uQżb�*��&���m`H`���<�g$C�@�M �k�����G^��e؁�$�9�/��L��L0�qCG!�(*%��U��v_�++>�೵{��!}ZR�__�O���J�i���s����I)f@2=�ji����I/�}LC�	������PA�dT6D���]�bUqi,=D���H��&Kd�&�֕�Dж��n���jP��]�3�ېD9m�-L*��[]��o�Ȗ��S�@�AVu������#����+�^:��j�&6��� �v�f�����Ĺ0喁1!�p�gr��/P�2�����n��_,R<�;�KV����_��"�sV�Go���$V�OT���H�5y���F�/��
�����j��_��& �����7{�F�a��a��B<���(�,�k��S2r���1+�<Rg���M���T�@p�I��j����G>a@�%�b�}a�¹�$�T�`�_�%fT�]�>��ڵ5ɕawc�{a�o��	.��V���������:�d�����T.�#�k5������.@v�q��ěj��L+TI�Z���S�`� ���&�"ڽ��y��p�?F��ЬԤ/��@����u��B�w���jK5�����ۂg2��Nd������jlP3����8u�y�sp�����Ѵ���v�s<c_S'���AC�G��]�ÁI�=��M�?*�a�_�Nǲ�Zm�;;%���(��fӠ�24�3�zn�Kw���"b�=��������X���a
HF����Δ�Ƶ����>�\�\4z��t�|Z�n�*�>�B�c��H�ѿ�ʯ��=Yܿ��ѶJ�W���>~ёf��E�c��,ʿ5���<K��׹�4��Y|B����6A��q�/o�GD���}4C�[Um�/ɜ
r|�R�٥<���W�;�W�nh���%�xS��@r��Vzk{��>�wȰ �E�~W����/(�/|5�ՕUM�Y�6ڷa�D'��|�C@�A��߯gB�nor ?Wa��5�6+ɀ�T�}&C���,4�dn�iߨ��Mى��k�|(��j{�%@i;��^�}t%��*N��AT瑎@"�pCMt�W����]�+�2�R��3E�����.p4��6ʃ��|Ͳ�qqp�s�̅�?I�0ő��*h�q������@u��$����W\����H&6��U�cx�I)q�fL�A�a��8�(�˒vz��fg���)���r���b�3g��y���2�X���ڮ�#oU>�G�>�������m�y���a2ѭ��+�����p��lt�e�KN��2#�����$��Hlc�֏��N2èt�ΈU<���=��|HN}WPs�?#&&U��5yN��T��$��b]��)Y����ׇ�
�9��%�L������������k��^�q���S4-�2�f,��
f��^�j�u��&�>
�r��٭<�߈�7:)�OWc?v��l�{G��h�K)��",�	��h��-݉�ޯ�|�V�����Ḭ���%�$�rs�Z���}M)�̺:��BY@gq8�0�����A��~_�5��z�	�Ѹ:y�1���p$tiȬ!+�bP���{�^;#{:������t�)~�Q5��+6Ƅ$��$Y~}�|B"�;�e�/�޵��L>��NcL��,|�>�(��v�^BJ�6D������wy�bp����m��>m���$8AJD"�sH�vwx���:l�nى�q.�.:�W�	����X����-�N�+x՞�����cʙ�(�k�m_2��A�6u#����\<P�D`����<�si4PR���d.fB҂������{�j��~q�D���B2�P���#�(XF|X3C2�X,�C�"�wL*�����ڟ�\�/�~�:��ɮ�2�0A�z��J�87u�06��/�3>d)��  ��XS������d����V�U���SG��;T�K#�)؁"���Q�� ��~�gRq�
�b���{�Yؾ��+J٧h�P������h�+ ��4��rj	�i#��,qtA���=�u�(�?t
sK� ��u��X�����%�g,�6��� �L�����##� ���ٻI��2��T���pJ�Ci[�fbj�:HFy�oGO+G[㉣A7	�kE�d
�͍��7�ǁ"F����9�o/O�wvh��F�hkw$033fM0����Ϳn��,)��6���i�6!��uX�m�J$lC�=hr��]�����y�'~����T-cj�d]?�e���3��DW����{~8U1��ۍ����+�]L�s^ơY�;=篸&r�Y�1�ҹD�ez̻��|m�s����~,$ۆg��<����4ݳr�1�w2��H��y��̝��>i�b�0)���q*<�N��[ U�.��>�I�R� ����0��RP_���
}d���5H��r��dM�a��nV�Չg�Ӻgk�E��������e'.1���R�.�i
D�͐������!����_u�Bg�&p���f�/�Q�A�B��4zCق/0v�%��C�5:�kpE�YƜwbE��W�E�e2�)�b*��(?���S)>Oټn�>���+rf$g�$8ي@�=~ӈ��GNj��W5\��b5�iU=�啕JuN�B�$���^ ����
�,}�拽�g8�b�Ǥ" _!RZ���i�f����X�܊����X�0k9�Vq��f߉�w����E��<4J�T�t�%U�H�^Q|�*�*�=�lE��%�����ؤ	��C�9�c�Wv���Dk|us�p��f��&Q� J���!��`"]��b@z�O����a��d� ?�Xz��zO���0v�T�n�C��a�}V�n����6F=L�8{D��nY�Q����-łf���j�p�h�|��XÀ�F�g݋A[`�x<**�u^�3A��αO�|��e�OL4_8�e(�fe�]�_�ڄ��u1��M�^��6�4ku.`Z<x�$d^D܅XK�l{蚬ybY��c�Q�Z�a� S̤bo'��j�����t\�Rn��VX!l6�����H��aD�u���o��Dnq���9����eRt��
�$���G�S���) hU�T�����d�}�]��!��+�S�[E%���Y��Q���;��n��l]���[�Y���<Ds��O\��vn@��3]��s�ŷJ�c�#eN�@�$��6�<m��-`���MQ��q��I�r|����͋~���m��,Mڴ��|�Ed�R�~(�R��]B��"�(nHr(D(�HQ���zSl4����k�M��W��q[v�|H��~�;H�fe}�.y�yJ2}�����3?
��(i�!�s-�y�c�8Ư�e�5���t.�To^ޢ?T�/L��3"�x\�F'��ܱ}> ����ǛN�捏`bAi��맪z\i����<�q��߮D6&�O��D+���]C�^�DP�yi7)o Խ�A����~ҷ�g�<&�����+8�Ȗ[k<V�������!�n����!���2���5!���[����>J2�6�
�e�i�*_�D�%+�����j�����)h���b➌"k���6���D�cc�\:��]�8��T����+�*RO> �^�&;�]<��'�e3����%9��5R������k��+:��$ܨ�?]W�{��X=��3P��l�@Y��}��A蒐�UZȦ����
P;�@�.9��ac�γ�\Ŀ�^ �+��u�~��6���	�Ĩ��gf�*���oЏ�6�b����@�)��>?u]^P%��0�kx8�o�u�θ^)Zw �����	d#�/I�'��z�0�h~�������f�>�s(��oΠ�Y�R��.�d�5�ͣ��gv�^�X�4��s9Y�y�d쫖�xB�^���n��W4��:Ɍ�J(�-+<|�~�HrOڑn�;�f��;�f��YcΞEA���-����x��9���H9S�"���T�k��q3�X�x�Hlg��ޘ�R�k��"7	����������p��<����٣]����yc�9�����#�� z&%�� ��j7��y��F�n!�4��ش��]�\����g�vߩ~%av!\�e��&�S.�]ԋk|#�R6�W����hMJ'���4I����i@-��=9}����&Ki��[����R��.O�:������6�`����"��XICz�Mm���x~�j�:7����� b�P�ɞ]�����G�j6a,����%c�|U�ͮw��s>��S�Ju��f��g:ѐ��\��X#~fABf���q5��Ȃf2^��Q��,�CBe6��KMcrn�!��
�=�u�C���n�msLH�ۨ�-��.�{{{)�$��V�ܨR�iJ���������$,\=�[^�i(<r೼NB�Uƹ�,��i�6#q«M��W���^�*�%� ��w؎�%��cŝ��iI��^Ø�d�^�j����\�����Vd�+5���'�����7�����3^�����k��ٞ�������1T8��`��r��nt~"�͐aR�E����:w�[�dD���N���hNϑ��ى6�*���O����0��`���G!��������
^����/�����=~�� ȹC<xCj���
IL�թ��d�%̍[���{U70:3���eߝ������8pﶸ#���Љ�p/�J6H
e�`�Ld��N	U��{��/�$�-��t�����gcu��:ϸ�Ylq��)΁�.=�XÎ��}d��O����2i�Uk�8��L��� ��tNȰ�V��i{!qS
�KPzX
hwI��!E5a�J{�aD�㴖��H�7qG��'����jVҹnt*v�"��~�Z�s�8�IR�LV�]�16�������mt���P�_�%��'�Q���l/��v�L�L5I��90H��l|iu�q.|����d�G��D	^f��;��{dgc����z�QL������n9�B�b �T
��ZK��� �N�����7`�֖$����5�rk�b�Q�ˑ�CO!��f�ǂ�ljFAk��^e�A�� �F�ĵs�3�+Is��F����5cX��חV�cJ�a��#��b���U�QdŰ��]F�A���,͎�hJ����Sf�a/�8�;��� ҟF��%�y�t��/����w��W��5�*��Y��|6�	6J%���L�4�QC7���m��QcGվ$�F`hN$@~�j���vEZJV�6�����qS9�98_�K��o��gKF���G��V�y�H�10�����A"_�_���:N����r�=e�����u>���!@���M��)�,�zP�ֈ�-L	�ڇz��B�N0�l&!�/_�Nxڏ�w�X^���slݫ�	e�Y��T{ަ�Qx��nM���k�:�{pg��h:���Refe@W2݈�Z�V�O^��ּ��a�G0U�t͊O����} ����83�Z�aͰ�tݤp��<ZV�
'4)}�<}D�z&"3%%t(�/�P���~~)V3���t����܀�uT\k�{��GR�aVh��f�4�%&r���>CT��:���9�ʽ���Й:m���Z��o��C�޸W�І��v��fc`�Ef�����Y"�`���U�w���P����7ͫd6��W����Di��t�&���Qͺh��fZ�����m�J�>@o4m��H�}�Z�3B���Ķ/�����Ck (Ώ�PA��Ood�&ȗI��:�Xy.�K��Á��ߥ����!5�D�3���	�ƛP�I� �K��	+�����X;D�	[V&!�>o��Ù�~���;[�K�R���>����ԏ��Y=p�p�ksmE"�<�zU���I~��+�,��㟒h��>�< �'�?w��1`23�\�V�/�K5%����
I��TQ�f���j�M'V�3Bm�Kq<���ݿ���q�p҈�n�k��a�y�V= ��OZΆ̂<����`L$�o�mژ�����:RKO�Ks�lK�å���`�F�4��,�7�O�����n������i��N�.�a&7��s��C*=h�o��l�����cc��r�h�*��C{��DL���{���"&��fojZ��?��U
|�`�8Dn�/_�A�j��PyB�<d����8����e�e�t�5��ywz8�t_�����*�4�g*�����;E��;�<gY�pb,��{��n��źn��}-z�I�tբ&���mVF�j0�:�?�y�2�H��$����
.a>a�L�'���1D���Zjf�5�E�|n��cb���r8I�؈Z�I©��`͙�5?4{?z2%ց������A��f�� �
��/p.=��{t��+�P�'`9��w�p���g�K��*zzK���,S�`��`8U�+iyI��d����c�p���ʢ�M���y8��O�̨mM�i~�����Y6֊�J)Q(���~V�$1���m�z53��yQK4�l�����O�<�iG�%�f.�z3ϋD��S�Ωf렇������>idU)��e�hKwex	�O���]��$�0�d�3���YW8�V(�~��5Ӝ����)�+X�]<AdYs�`b���3��`
�/�v8_"7�Oz��3�y5��1�
x5�T���Ϛ���+�d�b:/��zh�}�
�����B�|�m�=Y�Q麥�hϟxm��χ�:"�7dX!�uy�B	 w� ��DS`j���z4j��w-��%v%��ٔ��pj���M(<�b�o��L� 9V���à=��G:�o ������4N� �_,.��?%,���8�0���,L�Ř�J��, |8�d�k�j�雂��F"Z�@��k}�{a�=��j�l���Ɋ'��N&��Kx��ؓl�)F���x���IK<#q=�(�%]��7{@�ēF��'���+����P�˴�g?�<)�3d�տ���Z�/���q���jU��z�;��V�[<z �b�ֵ�m��9�U���;	[�WZ����K�T% ��c/�u��n�+#S4+:��%)��f6��p>�`��`�e�����/�/>���g?7�n�ۉ+a�:�{~p���W�#�x^�BȰ������e�Ϯ}���`��d���9�sHUe�m�0*�Bi+-q����)��
8���'��������J|�6W�BA�J4�hD�����:��cė���Gy����nN'i$����sDii��7b�%�ə ����OεVc��6d�/cS)G���Y���7b��7�7H-S�$�zo��0ye�EB�-����I�����f�nf?�F��W)��:;T2@��t���Mf2��E�ۗ�����U��'��5�n1�=�%��<�h��YVN�n��Z���v��rl�r�g+�v/!oҚ�"��~��\����0��X׹�'B�uƓ�B*��֩������d��z�މOD*���R%����L.8gy6�A���b�ܤ�����m�$�[�h)����L�P:�~�E����m����K�B	Lg�3'�{�gS���n���3[`��$S���/�a��[�'��b�ӼI��qJ���V��/dK�ۯ��t��86ku�>Z�*ց���"���@Y�B$��K3y%�I����Ζ�;�_�]���͸3���^ݴؠ�CL;Kc�0�nn��)q&V�_^0��G�#k�'�$,��y���}9J��?�<��I"<� m�ҫ���;��5'�Z�ГEP%頯TX�����>�H�,Cv_)"��2d����?�|NF�T'���l��Q��MDI�\�?��%d���|#���S�:��LT?~�@Z�}͡�	t�@��Z�&���҉3B�s��1�����{@�_�Oӓ-(�~�rW^���}(����Tl�#��\+]$�zrD4�rj��H�����C�ÿX�8��m)Ԯ�I�PRPȑ�|!���~�M�o�?�7�?�~���q���a��˩�� ���~��9��N/���8�Z�����Ip)^6n�U�v�����cf���(8�YEʪɑ�N�%���0�o�問XG'�!�+6�_Q����T��������5���H�1�W�):#�2`|�Č3$��ޥC�aR��hh<��۝��]�����i�ja�uiOlO��.��r�/ڝj��|R�H�S�F5�$S�L��C��g��W��M�o'��ϲ�l��Y2�k�$ݧ��xez�Y�
B�j�2:fu��&���l���
c>=����^y�O�uW/I��}$3طJ��AǺuĵȳ��=W�w�t��tH����sd�_�!���A�9�[]5Rᆥ�|��h`yI����Ss���f���m��G|�J�Ip#�6����oY��;Ư���e�棱�00R]
F��a�j!����U�GP�X���3�7L%�5�܊�ܪVjr����9���Z��V#S��o_J�-�u���o���0U���d^��,
2�������!�����I5j��m�^���J���U�[�-~x���2D��s�)$����5���B�rC�&nb�d�
�O�t �4@��vY��ھ�l�W��q~	��Y;z�l%�.��z�%|J	�FQ]��́�=0K���Չ!�8
��Jld�m��=_+�����b��D�P2���+G��qg�H���!LR���`,`��_kə ��K��U�I9C�#�F�%��8U������t����)j�c�Ȏx������������o4D ��&�@|�.���� UrQ�Y�G�c�C���~j�L#Ș�<�p	�_�=P!����� �p��s)T94D�5�}K� �}1�n�mH�fρp����YI%B5w�v\��;��(��jh�RIc2�9x3�TW��?g6��fu(1��v>��r�s��L���H;��X/}-�5�W}�Z G�u4g�T�E���(��}�Л3�r$�|c ��]�GuI�N�[�*�w+�bN˓�曂��"W�]3���+��}�ʏȓj�G'�`����;��̈5r@��R����vGM�'��S-;z$F{g(0���o�p�j�H2�#³3]AS�yBe�Q#C��t���%������V�S��9�T�l��is�5���6R����l�b�|H�����f���	�&��nc��$����L(TL �b.]BӠ���A���� ���4!;��ffH��^7� y�P�̝ҁD���طP%ՙ�� ��A��TV���&J!|�Mَ�(FAR���ӻ�����t�|n,�����M�~��4�,A1�ş!�#���i�,��Z_ɟDBm�G�f,.�Ѻ��؞wp ���'NG���<?�4�ff��zT��u%N��{`�LrH�T��4H?ra> �{�n�5��d!N�������b\+$�qr[��Ne������ȨDeP�� N&ko��n��TAk/Ӈ�[��!v�x�<{b;_| �旳>,i]��M{0V�ř����G�~�Q�s� gBZJtf�7�j! �Y��{dI!��H �`��1W���,�t���]�������C���ʰ�� ��r�8�5F]lE�j��N�Ӧ�E�_��D��ӏX��ƷˠI�*u�*F�N�H�E�|6M�<.d�K:�"䎅��v��s2e2������[��y���$�ߏ�?��skO(G���=�����D�b�r�Z���=?����l o�]�?�s_��N־l<r���l��/"�䩷��:��w�#��]ߐ|�%���j�\�~�@����+ݏ;N�,#t���
/��
�m���c�`ML]�x�8����s�׭�ωOr�����'j �M:�����#��@GҴ"��ea�bd�2����j�f�?�|�	\G�h"��*�Gn�<����<A
�����Y�N���mlr�h��� ��;�ײ>�7Zh
�#��"�G�(u$�?4&ԈWtRJ��I����ܺ�b�p:�#N�J�p��&�Dv2SE���S+3����{�2��c�5tN�w�y,�����R�&~S�4b�;�����(+���D�P���U���*�v��o�����$�zX�@���� &�F��ރ�0J��<)o����	��FH(o�a�ͽu�PF�Jr ��H��s<y�̈�C�t�l��'��Fj'!eXO5��D�p}/�j����7���������U�
nB/�	\�S�c#f tC�H����@Á�\�߫3u���8?�m2����V!���z�e��z��C2P���FȖ3��e��`��%�I��:�Y�X��S^v R� w���ZR/�x�0���t��刵�t��yI�~֢�zR�K����U�Z�0\)��*������!Î����Đ3���l\�7��PJ�����_^�݄q�$ei�S�O��)���q�#��p�Fk�һZ��S���@�D��Ƶ�C'Q�*�$�lp�Y�|��Sgm}pxKXlxV64EB    c726    1fa00������+��[�`펢�T���H"Jn�<}����/�'����׵3z�q�=t��D��H��jR�>�9�f�z��.�E�P���ݸ������պ���Ã�l�~����L�-�J�"��zY/��t�:�\�G0���;�j<0��v�h^�7g�O�4�5X��K���DzG�%	��W�4�V��NLˋ����x�qy��m!�Z%��4�J���<-�[�p��c\���u��40E8�}�GD;?�\��&���Mt����b��>vKt�ۺ��d�_4������s)�^>%��b";�����б�O��T$'�;Sb�=t#.	a�҈m�s̈́���đ��,�Q��|L �|���c�M�!���+��������t�t]�j
z�9�^N.
_���W�C�-B���|ճ��,a��	<�\�}�R��/�)`��������ZuiP-S��h�)�h5v�J�����Û�������8"*��Vì(��ꏰ���&�{!���C�=�6���]c���N��n�?nM�k�R��A0�7�Vm�1����f3�b�8��_D"��o~�j"G�u�}~:�S���������Zf�&�9��3w��{�qa�`���*B�R"��᪹u��e��j���c��S�`�Of�62`��z!4^9��x�'�XiǉM�8�_FFWT ^I���q���k����l9(@kT\_v��H�?���UqQ�m��c'�4��O�x�!<�Q �[C�ZIC;  ��ae�WH�7/]��� � �zwxv/*`DG�m ����56�4�]K79��o&�� �T�Ŷ=�9N]�N_�)\�c
0��c���M�Eg�M��=<J��4�l*
����\��l��Ș���~�5��MK���ɮ���wM#��C3�_��p>�]RΥnq�9���㈒��$2���b:Z�,MQ��N��;0^Zb)$�&�.��}��ތլ���%�G�pҟ��B�a��`�e,���o�.��ϕ�9����c� q��Y��ɸ-�{�Oڎ LUH�0���k�;�^e�����=S�䌮�XU+E�Ǐ�-#
�q�ZK�w�c9�v�J./���]����l��0�����ˏm)0k�[��C�"�� ~���4B>���v���0�N��+@�/%�J�7��u���%�g8��2�}�5����_�A��JH�m�D]�<����B&�qQI���F�}�t�
k%�����p����b^�	�����{iA�m���(��1���BhQ--*�g��]����A��=���኉Iq뿆c�^�29R !T9дe`��s
P){>m��!��TxM^ق�z�8xy~��+fB_`��.�k�V�x!�H2iï��-�}~o�i�U�|Xd~h?C��_g��e��GA���DG�}���{�=�؟��ġs�<���PF;���C7&Da#$��j(�H�B2N�Rq|����q��%[���I�!�1o;�����R�k�8ݕ�k�}5/F���OT�r����ۚ�upX_�72�pq�*����s��\�ꥴ��E+�H�u�芲���:�d���j���>���ev�n0I�^��ї(��o�2�bέ�'�su�5SQL�t��r!��
Hd !K��&�K�}0?�č=���*�E�5�R�0���#�:��2���9�h����Ui` !�_�x`���|����]%~y��+��9#,E����ͣ�<��ZsA�*��}ΩР��FE`���eҫ� f���i�t ���%�-�
v}SnU��8���1	q�@�&b��H�:\���!$�kjNFp���-Tx���S�Qgf'������4]�6?��i�j����փ}��L��|w��,���PHM��z�Q��;��o�}v�ơ�ۆc���zc�p(�_��l���b3T��{-0ۆ��9��W/�a$�{c��w�n[��-���E_���+²�EC����jZʿ h�|����z@��� ve����0��.��(U��E��w��T�SwO����x�~��<�H�)#g�
����ƿ0*��[��<�X827�o�����̛B���������K��[p��4�Ӿ6pZ%�@8n�� �^����\3!n�{��gF��)y���b���t�E�o�)!��_D7�US\�2�ͧ�I�-�H����#1K�Ink��38:pi��l�낶L.zn|�Gu�5��ex_�������N��X���S��2���L��!�!D[���I�<#KL�<��~�g���8�D�7�'�����A�zeWԇ�}틂�a4X�
v�3�6���(_$ؿ�����O՚7�Y�`"�S��9`���c�<å�R��)��U,ٞOa��O�����^|TR�X�j���1N�6}-Q7|��A{(�;44fݚ�d�0+����F�J4�/¼/�s��z}��=4T��Ң��u�-?+)V~6���h��u;Q�wH1��X�췽',���kf�D�k�����t��꼑4�`���n�v
ٮ��2e'���p�,��8wSk�{ċ0���:�N�-�vS��z4,����_��U �I�W�B���6ٖTs]#?;+,jeGԋ�<Q��v�=t��
��5E����Qq��s�kC
˵��}��I�jFr+����/x}�	�a�y��#��=���/��A��f�L7f���j���}�<ɫ���]�!����+�>X7��n�@Ȼ�{E0�R��KY�HG�m0�ơ?�����[p�����i�������K >ZasZ'�Ǹ�\�v�k�+�G5K�z�������gr��
^|�������驩L���LIQ �£���Gl�óWJ�h�������S�bE�q_1��P#5��?A7rW��2�?�BE��p�i�9�?�}�����0�����ź�J�f��Q{T���*)�J��y�C���=o/Tk3Ǆt���m̺�6���[*K�F��ō�ς9ΒѪ��|V��o8Vv1���>_��^{P<�w����<Ŵ��WRCT��;#fI��h�܅>�
�yu�sN9'9�8c�M��1� �-���Q�+N�������ŃO͔��E�<����`��	���u�\�̎�0.�r=��������ZHĂ��a�C�|���q����w3FMz9�M!�'�7�gw�e	���z�e
)	���f�N&C�s�n�ڲ��~mdOyLzO�S�&�}YB-��yD�e�;Eh��������wC4w�H_��4@	�i��6�On`�J��A79'M���w�JԼ$Q�D��?u� �=��$�c9�n�����c��^&=v}iwH1�*]�,�a?���t���Y�;�a���]�gě �����I'���zrU��v�3��'1�:��GQ���5�Nq�Gп-�����{�X��%�N��>��Xʅ~ ���)�sg����ރ ����z�{A=��'~m�q�=�����Y�q�ྭ�]��&
as�ǋ��Z� ŉO�(�/����ʀ'�zMX�+�̕���恞�\�ŉ:�n�?m\��E� ��n;w��ni0�����;�N�}���0A�".�p�]���j�|����t;�����a�&ʅA�ఢ(|!
Q�&��s�8������3@�\��	��aӹj	���jnx����؈�i�W��)!�]~�J:��W!݋�;^�j([�Fȧ$w�ʅ�T���u͘T:e0{?�4[��]�>xD�]>�0�����	J���2��/��A����,��(Ń����k�%����)�qR�k��nO8�5�B+Iyz]�}C�	_���R��i�n�]�L���8�X��W�{�a�����1b����h��Z��!k�_bK-���:þ�9���f���C1RTk<|�Q:Ϲ@;���R��y�(�Y�n���e��`X�NL�qS��:Ɖ���&��Wm�ʊ���V
���5��ȥ� R�,���R k�F�u1otc�}<�o��-���-$HV�J�(��C�[�ۧ�t��Y	���1��}\Ry��Bնŀʗ\�����S�m�9	9�9wa���7�F
���ܔ#���E�x�b�˰Whw��C5�qC{h!"���m te-���4a�E>�ϲ!�L�(�T5���$'�r��]0�]3,O�DZk��pO��N=*��`i�gMe���8�9�����,��L
"������!G�nU��J6U�A�w�C��%�}'��v�$���(��g�׊��jG�VI��#�k��k�����Ҍ�Vf@`�Ue�ŭH�� �L�xT�TJ�>�����\��)?�%�a�ϑ)��0r@�3.~FĆG愖��L9���-,�=��>�ᖈ�n/.����]�Y���+��9���8]��1�S���8d�~��md!�F�/#P�ױj}�F���� �F�Bu�2ƫҙ����Q!u���>��� ˺�BV��}��(c�g��i��8%7�۫U>��	������Ⱥ��˕���e�2�`��-��0ф�T�թ��e�e9WϠh6�k�~xyL�}D�H���q(�q$r{v�~���KO�>���M�I�ߧ^:�/���lYs��@o��K��1'�ǣ��H��?j<����*x���]�U�!mK�H_�=K�W	ax������C��Kz�Eti�����������W��'A�{#�O����j
B������V�c˗X�����.�85�����r�_J�rSC�#d��#9��@/IH�'	����[�01ܦ���Q��R�4�.��
�믭��ǉSa��dW�cd;z3�����<�����/��̏{�f@Cd��O�y6�k���BM^���t#jRW:v	��y�8!h�uS�쐰���ٿ��[9��R��I�5��@�e]`��ME��PZ�4[I��2�X��'忪�t�W������E������a�D��������:��� �P�'��C�� �%�öӖt��@s�kϯ���a4R��]L�b��6-�B�b $�"sk���[.^aJ��p�IT���¥��dþq3��b3'o�4k�#6�4�#���	�NQlAx�H]���%�A�TSF�z���$z��8�@��k�m$�#D�/ �w�n�U���t}VD&�B���#��;���q�\�q�S��g.�m*f�̘K{�!S���Wk'0�7�+�2Icǖ�!�Ÿt����K��ٜ��@�Ik�bh����k�	ō:���^Wɕ�@R8�9J���8�($F����6bd)t�-��^ھ!T�+�IC�G\�S��}7^XS���4�$�P�z�e��Tz�5q�I�opPRɁn����~�g��)"��ɠJ�k�n������a�Ң�
�*���#(����A�d7o�_����Ej�ћ%���6�"zf�=1u,+�	�k�q}��s	ҪK1<-�[<;�}�����ªh��IZ�db�>o9&�%��6�B��
1�փ�'%)�F��A*[�����R�;qo�/5*y��w�2���5V�C�T�p��G��)���u���2�G5����$h��1Ƹ,�&&cf�l����"��� ����*Kઘ��GFT�/����RLZ9Z�L�Ü�뎘��̈́0�@w���?������<�N�T��X����~c�3`Wz�n���h�����X���>请��"n�2��Y���BT�k�5qt�&h�C:�/M��!�.�M̀��i��HUz���7Ly�Sƿ��˥��OIv¬�8��|���,�u��iJH>�Gн�󏭼@�g����?�Z�������C+S�HWFϷL�g-=�.����/v����r6�=FrV{tLf�9���٢���ehȞ�����(j��-X��-��~�bȃ����i��4a&���M�U|��!��RxF���P�j1��Jx$����*����vsےU��5�}��)e���L�lǮ�������}��2���+~|��K�b��j�1# �ʽ~�z�4�S"�4�����jѮ}��a-V����7,69��.�w��~����>�zW�Dm���GZz���[�~���Vc� �z�zܤݒRG��� |���:(��Q�'$ZC_ 0��?3����0&[|�*��>g=�3�w�6�q��\���V���Q܄}R���j���%c`���o�Tᦲ��%�'�Ê%�:FK�l������Q���Ơ� 6F���7d�+&���lڑ緒n�F�_SL|�����rS��_��	�9Hʚ$i��ف�ǔu�pwp�;fR9ޡaO���oQg��Ϳ�t�w/teI\]�_Gb�G����ε�"Uy��d�s�d��ķ����S���@y���~��)C*�j�Z�`;��CY�NZ�s�ǝQ$ ��[�B_0ei���웹�4��~aVG�*@�ӎhU���
�V��6�h*��!سu���_A_��'w�� r�g�k9���K���� ���f�\xI��@k�kj�)`����40o(�ѩ�ݶdi�� aP�2�ϠY�ޠd6�F�N^2�8��*t]��Ի�[I�J�p[�Cz&*�1��]Il�J-��/uQ���>��,��P�ܩ�<2�/$\�3�\��n̔bl ���J+Ck�l=�&��@0�c�d�Ʋ/��Q�(��_O�1�:i�,����-K�%���\SR���{�[�WA\OW��Sts���G~�H5$ձڛ��Z[�E6��W �~����g��T��s9��I���]8ދb8�ᇻ���ވ. u\5�C��u�%���D+�Qs'O'$�K%���!b,�'A~,�ay#�%�q�F�MrWwy}�����r��ӄ(=�0����� �]��+��=o�讶�M@E�-Lx�4xf�7�?�V]���S5S:%�(�;ɣ�,���s�Z@�.�+��s���}o����\��$5 s��/3Wn��Qr�پ���K������cl�`o��*JE?�OVb��D�Ǫ���{NR rn�<L6�1�;�I����{�R ~����+��5��6�!�%�b���eH����X�K�M�:0�ܤ�u����=l��$	����jai.�'�-�َ�r�
�+>���KOk|�&W&w�X)F�Ն��{,�~߈Z74�G����/Íc�
�����D�4�м�ɓ��ߐD�fR~�?��σ>�I��@�|U�'�ʙRH���7��&E`Y9G�wc^(2��u��70Æk�	 (Y\��gaGҕ��ө��/��WF�҇Ⱦ���ךۙ����*�>C���HR&��K��|H��ɓ�d�$ �]�ZI�p~�e��*&Տ�n�����=|ʆ�� �D �+��/�H�ҙ,�Yl�}VyOU�4�B)����RG{ �Zل�?ٵu�(U��T�]�۳�Y{)嘝�����a�J�:?���!JDpL\L�1{M8��l�O�H)'��\~�?�<Mvt��#P���~��:�"o�ȋ�vL��Zyﺕ�{~�.�~���5Dq�h��U��M�=����	<��hhFU&b$a���:�5�W�-D�`.[0��_�=�!�9�h1y��"�p$ܸG8���ؕ���Qu�>�;�Y{rYF���b�3a��$�q�X�Q���Vc�`"AO��]�p���:�'[���VK"�`@��8��͝ ��8aE���6H���1��=�H�^PV1r��>�Ҵu"�e`���'g�cHL�*�D`�'a�0��a�/]L�ıR����8�op���[	��B�t	���3�M�IJ͜�������R^_"ܿA��}l�*xkP��Ns	)�O��h!Sg�å������}-��!	c��q�4����qE��@1�yRnkLhM�6��6�����.H��m	�X9��4