XlxV64EB    3a3a     ff0�i	,�2��[t쪓y�:�g�q�T�s\Ol��P՗��9�,�b���<[��Q~ʱܷ0�f���N(..�n`E )l;HmYO�����T׵�ɏ�����(�n1.{B�@t�����a�+���8�G���%K}�utҧ�?�D�c��U��[�$N��"ֈ�v1Q%Tîm�Ϭ5{!W�A_�s%O�lv�PH��:Y�/�C�9,��].h8]��ƽ@�yJ�KS��f}��y�/z[�ϻT#�
1%��$_/�\ll�;?�~LH�i���v��z��σ`����M�@�{�	��Tƾ%c�26 b�P�d�sY�a#x��L|F�$������/9�p�vg�}��BOW�� �H���4FCp����_�<ޟ�#�4ܘ���/'�A�����)��o ,pt��E�х���(��M���k�u?�W3#���4�c�>j��,����C�g�
��~��v0�6�s��lw��(�O�>M�뼑e$ ���U�������T�\=趉��:=H��\��d����El��K����(�+�/ɵI2�(~��Tx5A���Ë�6l��7و}*뒻=ED �p,A�F\�gs�X�o���1���5�^��E����3
!C�$$�M�a�aۜVC��f:X�<�1X��F;��dQkp-z�-2�Ɛ��]s�H��'��?
D`�]V�m����evA���7��`��Ã������`u��'8�Gŏ��I�Pl_��^�������O�4��\^F6��*���o#��M������Pv::T�aF�Yx� �S	����!70^��)M$d�|V�"9��US�{��Kmb�N�O�B)���r�����#xb�|�R�Q:b�H��:���6�d�%�H�����ݼӿk���C�3�&G��,����UP��|�^`��r���,���؈�����3K-l;|w �����xtN���[2МMe[r��"k�(���|,������?��ef�l���m>�c*���06��Y��IfKn8���3�ao�p���$�w�Fro�t1B�&Y#��A��y�M�h7-­y>/7��Pg�)�=�NZ=������_���6޻IL�26��i���|�X&�`�F^p��a�7b���_��:���]�E=�'�|�|��R�[Y}\)5L�T�>#�]�adMm��/���gg��ZKSl蛛�A��.s'��r�O�O�,lh���(	s���p�Yf@-Еh?/�VS�-��QA���Y�}4ȉ�O<�ޓ�������s�l�{"J20� �%�"1���I���6���k�1��E=��w1.�R��L�E��+����c����Gl_`i��vw�o<��I�b?!7�CS�v�"�ء�[��VJĹɬ�y7�%7j�&�`�:�ٽ�=�?���[��Rl!���H��"��7pr�#�M�>M^�m���7���7:|pp����p�<�1����W�?SI��y[���\���5 L�9�.o�����T�l���/[�6��6�U$2�9~�	��`���C��r1V������n���Fշk�I���,_���P9B���k�X�F*Sł!���+~e�o�
 �*�,E� �=�`�"]��=���J,� j������
D~6�����r4���竘S�BG��@Q�D@~i���tE���J�p���͡$�� c]1���I�$[<��A�b��/�լD��U����C-t4���h�g����JN�c�`�ݗ��6-��	����`�$��� ��e$>YP���-x��˯��-"����~��[�ꭦ���8�+�W]OQ�6:�����7y��@/�{���,����?V�f9�!2An�����2�������kC<�__z�Ns���	S\���v�������>��_������I�ʀ��(SP7���(����Q]u��0��YW�fD+or�ꄣ3 l���֥��P%W��л�#����콧�m]�4�/F �U�"2�"��k��yZ�j�#N��c��'v�Zɨ�qaǧ��l�s���0��� Q�v!�G�0S��M>a�#�2��%veQ�y��{��ńj�$���U�)�ƕfyu(�ti�mp�.���-4)��쬱���gܰ�"3Ի	�F_e�,iDh���K"�)�%�\�ܙA"�# �����Oo�K�Nr)+W��^`��/�V�2���w�6K6JvQ20��}Ab6�jh1Rrѹ��<�.�+��s��G$����'���CZ�]�7����k�KjR��*k��*�CB%t��F8.��b�X�R�E7�&�H��u9����øx���h{���PjT Z(��3
�5�Gj����{gR'^�jN[�Zh������y�0�i���M�5 Nf�V�Ltl�T~�s/�% �o��q�Ԯ+�q0Zm��g�m�>�gyk��v�8�7���D�/��J��<��R�����d�O�䪹�u�Y��,:':2[����=��s[O��״����cYz>Ȋ>����V� �E�ў�r,�����o�%�M`��?''��Y��g ?�I�[2{�������8�;�8���_�	���	�usئ<0�Z����<��T��_�f�G�3)���JmJ+���F��{2�ļ0����=7�2�x^��GA�c(�΋d�v�ޮ4*F�x���p]ۖ(���X����A�h����� ��a�\	xѪ��!C���<}-f��H7���}"V�䟝���A�l�m^��)C�^;�=2Fڐ���!�~k����X�Ƶ7�������CO+�5�C�i@�>%4����0� 7���w��x���;k6�����s��2/8C�/�q?�Y��{�x����J�Pu��ǟ��o�7������j���"����vNʢb���w��?G���m|z-9�Y�6p��jtNhET_�g��"�.�>7\.F j␑���/�p���si�O�q�i�9���^2x�=���Rz�<���@=���͘����M6	�m�勷&ҵ��� ��&������>���}�b��̨�����n=�³�%r#�\]�d���+����P9tw��v���h�k�:"o�݉�n��~��.��Y�:௴%�ޘ�|���&w��\�n��+�M���PD����R��m���J���0&����Q w�,��MR�U풂E�����!�#�������+�q�-D?VW��0���Q���5D�e�_�%j�:	m5s�H8X״N�: ���JN�,/�_ӽq�`�d��ӣyR�x�Z���J��P!jn�KQ�r�ptXQ9̀�̼:1�[_�� pǢ,�	��lY��~
�gX\ ��	��	���b��y(�W?^q�Y�j��x�^��a��zզ��8ig��Ԏ���oK��ϥV����f��� ����!���8���IJ�j�z���qj�Ig��,q\�0$���y�l<��L\����K�7���T|Ѝ�aMJ����]�4SbD]X"7\��Oǆ"�,�4):ֻDe/)_Y�ZT��5��`�=QY�V�Dd$�vN���;L9�"�5��Lg�`},�^O臯��v��;P����*YpTH���39v;G�o�	�i��ΕG�����(ad=!�|E�lF��~���B]0�T��CND����18\��9�4���Y����$�U3�~�E��4y۽U�E,��h}r�
�r����W"&%�amyu�-|�"�7����ta�>w�� ,�B�}�� ��4O��M��1�aֳ��׺�n�h����1���-�]���(�Cy������ۈ����U��޾ef$n��uQ��L�{�Z1��6�����o���[aO�+�cW˷o���ߺ����k�&S ?�����W��]��Xa�����eיQ�aɗ��6��+����z�]y� X��K��A{���3��"P]4��@��