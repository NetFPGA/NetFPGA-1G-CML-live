XlxV64EB    1846     880�S����"�+vA�rw-	�2I���~>�����QШD�%QVFvۅfz��U�D|���e�/�&�L��}�~FǸ=c�c��2��T���v��#x#-�h��sc:��/������������޼��tr�I�5�3RvDWg�����&��t02�W��H&n���%^.��T�9�Wκ�S�C�v����}_ f-̈́��������`a�������jܰ5ђ���b�8���.�K�a�}K5=(s=y�b��uV}�3[Z� iy�4��J�ZĻ�Ș'����I���.��%��� bО2�Ap��p�=jw�Q)��0LR{B�ϼ��;����b���rQ�Ȭ�zۜ����ݱ^�l��n�|5f�b�>J���pJu3yZ}�,?My�*v�"�^G��1����(�q��L�K��J�j�$h��Z^�7]�`}�q�
��bq8�V��Ik�Bߪ�(>�M���\�a�r���BA<\|������N��{��F<��6!;h��o��P��������i��ّ��i��"C�ܟ���ö�"���D��R�e�J����*\�����~�a��;�+;:�u[t�=4��ZKR���v�?��F�:.䍭��'�ڎZ����ޭ"��JY.�-���[��I�(ڧ�x*PW9�@��"���qp��Gt��F��k�ďyo<���"`o0$��]êH�A	}\Q)Ł�wŌF9L�??�c�<v���
)���3u��	;}]��H �}�G�fᰟ���q��_�Mt�۽dQ<�BwA�a��R�� �v��{R.����s��.T�����b�K��n���qqt"�'0��Ya=�i̓[*�q�Ђ����Y�\��h�b1�롲�b.�,�+���UZ�L�=d��581����%�B���++����S���`��4o4�����-��$к�#5�@c9���^��%�[�qx`RI8e�a,�^����_X&���KF%��W�E[�y��}�%K�J�.��f��_��I����7ht�s�#Ι�2�-W?�����ھ���~m}d�!/!��e��B���Z�]1��pvG�$��ˏ.�\PL�R���t����Op&i�f^0Ѡ�� ��2�z�>g���+�KK�D�u���NBrqp	��2hH�1��X�_Mw���N�f	:�,���r�׸.@�M|ytR-W+�P��s��� ��c��7׬��|yW�ɓlF�t@�~��O[�w]=��ȼ�%��k�+�)&.����L'\��e\\�,Ȭ6��,f�H�Z0ѭ�����'��`�G``�Y	e�¹'�]�jy<C�8�}�)���<�)���(�e&x�O�-UE����j��u��-x!]uǥG�'�q�l�A��K�wڎ!��[/�io�1H�1�6��x�_�>G�qa$4HXnh��߲���$�K�7���X��,t�9/V35�0L���C���x	�����劄��, ����;oZ`���.\���=�����I�b+Q�Qh[�v�H�1�[���pP'4VqgǗЯ@���@���`8-T�5䫖 V.ܰ��ʇи��� J�/Un7;~k�N�̓k������E��+l�sG��V���K:��KڲiI�����g�K	��.oD��q�~��N5����	�z=� �b#+�V
�X��Y�zy��ͯ���)�KƱoB�����]�\�_P�����Zk�x��2�d�/W��6~ѯU�xc�C����yLgM�΂�&%9��Qp�6�(A�ј$Tn@6��?wC/)�{�)I7`ih�cC�-1����i�@2������vuCY��HpcQAu������m� �c줏6W�\�h�_��-���,�'b+b#���l��3P��tԴ���M�%�'?����-�R/9u:��q%�]8~4�|:��]��ւK�;��Y�:�S8蚣��a�ʁt���}��k��1�y��:%����q���܃��JuÌ��1��X9�����ϯ�DMu�Y�����_�"M
fْ�~��h9O6 Qw�jf�R���j�(�T$$W�0΀��BW�<��� ��c�$Jʘx��2)n�C# 5r ��i?�,c���c���������i��ޒ�K�J�u=3���ҝ�