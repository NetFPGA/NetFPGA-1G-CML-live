XlxV64EB    25ee     bd0!�!<=��f��S��(�d�A�b�vc����I'������$�)�5�YtP�Oŷ���֘ ��a^���K0��<�M	���'G��(XXFe���,�� �X�9u�a�gf���n}����@���F0!	P�
(�>k�&U���{>kS���!�CZ���hn�0����,Ư=���ճ��:� �.���M�+�Ħ�˥1���b�b��櫙��q<T�<o?+ zY���k�UMT��!�̌�g�ES�����F|��R�0�;t�#p�~�"ES!��F�x�#(�rq�aLn�����O4���=��#���vY�2c���8!���"���h�2M������'k`D ],H���쩩�*; 4�Vf��%"�P��׫fx�/�U��wF�����LL��M ���UuV�c�V�{��Z�S.Y%�0������Q�qhŃ�3����+�2��<��iq�HЖ�P�ܻ����"-
�](T�^�+�8Z��i0�[s����D�8x�ݑ&vM�S.Կ��z�"���^�P�^M����?_��hQ�< 8H�#��͉�����a�e=n�v~���}���m�t!�9p�hS�~1�F�\̯%�2R]Dٴ����/����B��
o��d��m�6=�Ғ�u���~vK\A%1KBe�C#�qqb� PʨY[�Z����rn;C���y	�A��BB [��TWy��Gj��D�d���x�y��p�8�AI��<�?�qJzJ��H&[;�������05�9͸�:S�=8�rS$�y����#���&�A�jjaXt!E�a9]M��uT��d�$m��L��:�u�;��	�V)p��פ 1�ʷE���̆DL�����$^N�ԝP��g�ik�����R�,��S~8��{>���҄�"yNx�Z�������2��;���aLfm�E "m������ۍAޢ���շC�1���w�E�"�O �\����T�/��r��n[�#�"��Rqygw�dء�49�rˮ6��Qs�L����v6�Zk�+�/��9�6]�:��p����#w9EeEF���<$���ͫq�e�*�@9fiyZXh[A�,h=�8�P�^��@[-D�!U�H��㾍�����D$�Yf��	�S�T�T[�y�����W\\u�{�x���e��\���c�����*�L�	z��ە�V�	f;䦂�f#�5~���P�������ǟ��~m(E�[��[U�W`k��o����[wP��4ҜR�Q����B�Y����:��Mg�nV��,W�_5\.�"ŵX�*^�V��fuA�Mg��.��Uy�l����17��m���Bn9w7_��k^�x���w.�5x��R�~�2oq����Mg��&x�+v2��	�}A�m�O�-v����b�ia����1��tǲEi)�O�\!ƥ��%*�$ֳ�eP�6M%�7�#@�^.�w�k��A�WZ�.C�ےC9�X?L����h���~4�T���%��J}�XbK���[�3�E�[�BұӉ���܏�}�{S�N�w�8�Bui�7֠�z�صU�Ac�:)bm�h(�LV�;�U����,�|Z�����X���g<�`�U5����$�]���9[^͠�  �"�K�'�����YGQ%#�'ִ�لyDt��X� ��/<�������e!Shq�5j��=
��ݹ�U�0���Ր{�fj_^z�����q�C\׆tW�G��<��_�bePyM��8����J����b'6)�����j�"\�����_tRrS�<R��L�f��a���T,\p?����"�q�%��tF�N�6�L���E?_�_����_�4�fg�B��5
�r"s�TgJ\�!�sh>�^�4�~Fm�N��3��K��\��#�R�6N��Cտ��15�fV��we���V�&#+�=Ng��y�>�M�vD�;��,t�.YF9/া^� 8PP�`�*e���1�{��<i ˌĿs���<4A]p��f<{�T"�7u��<�΂��X�tu<Y�nQ�{zl�_�h���w��銋��"~{���W
��O�L�����1�J(���s'3$�Q�����B��� ��u�:V��Ź�qL|�3-�@	�8�;���H���yf����/��ϰM�B5GÞ��G<�n�N� *�Z=���訆d��(Vް�k�q9v�Q� ��d���9�W��)��!)㨈�����'��}>b�����,�j�� ă���_�eT�m��s5r+22+y�~z{�/<EL���v��%)�4��#����2n��B��u� �-�����0spTevV���M�eЁ/h����{mr��If�'=�c��d���:���3�����h�oZ��	'�9�js�&W&(^����I&��m�u�H��5˶Щ؎�oq�|��֧���h�d�t� ���m�r<uyX�H>AhF>Fw�r�I�M%�\�%;��H͘�
䡝��qH��aV�S�V����;`T��^�2=��ʧl� �SF6�$Q��!.��.
��Z�L��dY�5����@�*��3B�W\��;�0w�m�;x��s=$~D`��i�������P�׬�	��h4��y�;a,�cq5pl�l?$���5�m��+���[��ꓠ=��?G
Z�gN
ٟ6����HT���:�1�Z��za�-������M$��	4��B5�	";�=
�/	�N�0����d�4��ּ��5:�r3v��Ei��5}�~Ǧ��R�m1+*,�zյ
�cM8"�0	�~q�O�����T��m$6'�
��[��+�mG���4�`H�\��������?Z8������Ӄ�]�u�	
���nE� �zg��0������6���x�����2�]�9����g�e�諾�:I������R��ce�_��  ���fa��.��*A�k`����