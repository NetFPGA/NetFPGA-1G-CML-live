XlxV64EB    1928     9b0����n
ղ�Z���a�t��Q ���#�P%�!>��������.����R��i����7ıcblz�z�djjz��U!w�1�߄��p�9��o�m��I���6۪ȳ��標;�
k����y��l���_���ԙNǩ��:������37�������v�wL�c��Kfb|^�D�<{"���ax��OV������<3E7a��2���u~��U�7m��Aۃ�v!*��^g̜�9�?��\��,PH{0R�] ũk,�j`���"H����S��j�1��Y�����&�(�E�
���Ε���<��W�D2M��k��{ MB�#)+:8m��x�Ez?���]�#k��~�r���BC���}q��N�#��++l��mvL�Q�Y�R�4�w��X.��%�'5��,���e�*k��U�B��4��p�� ������ki�5Pk���j�~��L��?��)���K����6�p�N,5<�zc`B@s�a�IK�<0T�`A��"�IO
����� ��pp�]Ur�`X�M2Pe@��B���%���������=�P=�&�jaL�&&���\�뮚��5�ܹw卻r�V����
:��;-Y�
�vޕ�O���Q�<�{u�;	ǯKi(@4����'QG��i��=���_����,XBU��[���!�b��
�*'�Iǈ��p�U��Zh^�zg8m��|tO�M�M�	`�?)�K"�~����S��,X��K������FE�*��&�斈t��e�޺�g�M@/0!��|�Y C4��.���4<��c�����������_m5��F�o~�R�y}����鴵-du;g7��Dݓ|�Ǎ[�n�F	j\��])C��u#�]X}����Ԫ�bU"1�D��-�=f"5�-��X����J��Z�W���d�a$k���/����ih���������ߗ��M~��'�����<�d0=���>�^iDS��X�2qI���6�zB���HxvQH��V�/��CS�EѤ� :{[���|����7##ڄ���fQث^�, 8a�r��kK�O2�w�N�b~��^<oX���峵�I�����B� �"?����/���%�g�`b'�]
����`0��\{R2Gw��MZ0{d:�-�i����e�n]{��;�N+����u��q4%{�����i��m�#��d����I�߂����p6��db��p������Հ,�	!6�����RA~R�i��<=^��/�BlD\(�!2\�LJi	�%�!�$W��u���~3��ㅋ��/	�*_�~"�2q�����9�J�4�
��l�R�6o��
��e<�ƭ�@�ch%U�<!�BJ�:����t�4{s���{��e�<%&�s�n�,NͦD�c��7��y�]��~���WiSÍ��{D����v�|!̌\W,��&艦��a�?�Q��*6�$�Cb��l=@�p�S�\1龔H�N����;��{��f�Ӌ�G��TK�*�<>���U�W��W�:�bS�~�h�G�t�'GQ�8�P��7����~g��f;��, Fg�Q���1�D.�v-�+�Dz�u��3�eo�ĔN�=�lC��lĈ!3.� %��ǡ�A����Lf���`d�@M;C=3%
 �����}LS.��k�r4G��F�<�$�Ʉ�ٝ �q�܏��M(�<��5�M7E��絯&��;���Cw�!�
�H���i�Vև�b��(�5ٟ:��B�!@/����~(�M'���%�)`g�>��3 �f��[��s�%E�,q� N�2�S�k�Ƨ�3�*�q!��R�Y��H����OZ��C�E��fI���=����2��'�t�>�8�n�E.�?̲���L�Ȩ3�q��6�D	�W5��	�!7/B� $�a�b!�G�UsW���le�=Z�f�x��av#�ʅ��ȟ@O�j��V��}ٽ]����|;�o��\PHOe�^,�h��p�
��J�/gzS�"�A��K��
�ev���=�"̨��h��f�����3�������N k,����4�{�Bޕ�u�A{$g�1�k0F��"�J?ƅ!��?ei�1�Iۚ�T62_2*M4��m�L	$*��cڢ��@��/k�ꁫ�պ?�e�?��3���^~ya�Ȩu9��Tү�v��qdZ����2z�K~����J2���G��v:���3F�YL��լ4a�r�����K��C�d��YnZ��e����I�ckr@ֵ��,���9������T�~*hv���T�`9��ӳ� iC�.����]i�C(Qs ���w�x��G�c��鏉�*�Q��:�:u��Ҩz��E����'�?�����&=ӧ�&�ŗ
;�~k-��A�K���W�u�ŧ2{����L�.�H��t��ʺh���Z�f�>,���B5S��M�ϊ��