XlxV64EB    fa00    2f506��}r<�t�L��mY��!�K�K
	!��48$%��H�o��DK8V���t,����z��2��˒�'��6����\(��Y�n�l�{�dj�S���E��u��ԕm���6B)�
�|�4�`�̣���h�l[Z�FWp��3<���|��(��'�xL���N3LA���|�`���{�Iy�I�k�m�i�ܩ�JT���zB�(��l��X�떏 ��5����W��v���5$���X\��*W�n[��uj�\����_3�G���˂I>$߽V*��̙�Sb���S�N(��v�����r������^���rң�[�]I߶u�J�]�e��1�
�1B�A$���������V����k�6Fj�������]��nK���}o<��N��Q��m�_]�0���f�hH�f�;ct�gK�w��`VVY��Q�f�0�EQ�DV-���`x>Q�en�jM����9��S�k%�4�Q 1ɒ�#Ѓ/�a��S��A�����H�����U���5���������}���A7LFUV�!�ي�<��[���E�Cx���j:���-ڤ���3&2�*�M��w�-���Hf��Z{���zzF�f��э>�[���UL	��V�1��z$)0��Nu�t�a�	�dֱ����O��v�Ҟ�[ٹ(�uG�:�(�`@\��]R���t��N<S��
�(AD����3��.������v@��[������;Ө�md>_,�����D|�.$�0H ��V�E���E�;�;g�{��{�N��-*M#!	yL��h��b��W��3{�3�	 z#Q�]�$:?�/��C�|A5�b��>*�1s�b[��`-��g �j؜�R����~���R��Q�Q= 2���>���"�'Y%�څ�~��(T,V]� uՠ:E�sUς�I���.��i�j�C:Bw��{䊨�<�>�n�͇�p����v���O�O��s�h�d�&~���L@�u3�V���5C��PQ�Y��z���	�{=����8їD�k�p|�2\�$�[7�!Z���ں�j/]����Ӂ�:s�D�rC��AM3j��=��RY��Yy�:T��@64�Ε�aݔ-��b���jSuåJ9Ѳk`�����KJ��g�=HG��
_�>��vr�]='*w���*����&~NY�Eչh��y�P�:=�&�k�u1U���[�U�ɠ�UXv�l'60q����¬�u��k�H<���I�.�R6�k�\��e-�+��3�k�"��������2�*/������U�ܵ�xĜDu[��1П覷e/��Z�d,����{�5\.XI�� �a��kL�|5~�؆�奐�q���E%�-�,\as�,�&�!0m��P2�`���$ asyik��W�Q؛ĬH�l��we�p�Ą]y�i'bM�w�к�Yb|�$v�PT�7�Rn�CJ�6��_�3����%��;�)VQBU����7G �A����8��t��#}�g��� ��Ʀ��zl>wz>�P����,�R铢izҺ0�G������h�ڃ��䪭ʚWl���{���X$Cb��S�FUqF�\i�O�o������ȩ&@�yۊ7�h��鷝��8Du�1I�T�Ȅ3�M��T��4b���"��3(�eO���g�����xK_Wa)���vy֝C{g��z�3����.�bŖ��1e�ͽ�,j�B��﷛�Lg�a$�4^�G�]��!���Fi�c�����]
��6�������}�m_��mՉJ�A��P\)rd?;�h��WL2�nت*�3�r֡	�*�˰���A���~�����gs�!��F{̒�ab`�p%m*�gxo���H��^nk܄��t�:0kh�O���C<���:�i2�RZ�m��df���4g�G�
fH�bb���L�����.\P.��c81��#@*z���Ņ�e9juJ��k^XYb�`G��U/�m�d^��sZYԳ�<��1޳(��3�B�W-�WK�q�����u��'���=�UwbY�z��2L]�y%��g$?TyT�7m�	�w@yZ!�Еq���n�������a�/�+&���ȗ��ņ|sx�c�P �������а|#�<��5�����tq/)�e�8��8��-xUGSϓ�џ��R�g����ϭ�SGJ�MpTĽ4۰�����dyj�����[0�)��NU�5�򠔘�����"�OIJ�D�O%�&��b�Qz|e�NގU���r��pE���Ix���6Tթ��� �or�Y���,ղ�i���m��؂��S�f�r_����P�*�8L�Q��)�J��Ǣ�Kh��A��3����^�,�ߠ%0�m^��Z3�"�hG.b��{Z�b5@�B"��ݶ�;�@��:�����B��2:�G�-NKɿ�sd�ֻ8��2�k	R#��� �jO�t�l�c�E��hy��0H�솱��4���D)o�#A����K_H��W+J]�́4ࡳ��Xk~̣����DkY��v-:�	�J�Q��7����x�n&�^wzz�a+N��GdO��uVnk+ؒ��ə�]^Tl��ִ�Q�O� �` z��$xLn�c_S��sš��-2��V��%��Nq`��1c�
���M�8g�E�#��@Pΰ��Ӻ~�CI�Y!�9З�w�Xկ1��A�}�A�>=�2��[�[���A!�Ѹ,X0ǥ���Z^�^?ݦ�%>�ު��zT8�0+�놋�Z�z��Mn�i=k����\�"�d���Sͦ�)�t�[0�#��D8׽�qA�'��!��%�����|:kQ��2� �u[������U��bY ��|¢�L,��l��g�t)� �+*�C�WM�cD�M�����B+�r���҂q/�,�0Z�8��9~����2q.�J������Jf��
,.��Y�J���6��h:��?8�p�[�j����Ǡ������Ü
�Er�I���"���_IR��؊؉\�D)^|w"bI�N���"��@h��+�����M&�x�ߟ�������{����Z�S]����.̤�a��]|���O�ոq4}��flq����� aE���\C��&r�9��C�����s�dǰ�aeo/�~�V�Z�c�R�ߨ���Ed���ʦk���N�m�>7��V�x6i��nm��x�Z5�8L���.,��vCaI��[M�qխ|���g;Y�1��r_L܁<5�Z�Ek���L���"N��L[� -���Q�ȩ�ggBX�W����&9��o|�#l2�`�{r=7�l܊�=�ބZ�����+i䔵�����5��u���,*��´�t�;5 Z��_X��$ ����J���xӪ+�L��W�-v�ύ͕�Y�$����&�-��aW�I��X����e��A����8'����x��D݈��9��w;��d���0�]�G��O+^�[>T(4��-������q�~䋡"�84[H4�9~�1�Ū �B�$BS�2 �2�Io'���h�����s�d|�H1�m����Z=�UO+����z�؈g�<N"w ���T`�y���Æ���o`���ZRS���g1�X��?�$|MU��m����E�^g���3�M�������E�a��eq��8�DPň��u��%���[Pϓ�?)�$�"d��o���&�ϲ�F��f�	Y��n���1��c�-��_��U�Z�I18�"軈��̾ϝB"i�1�
����X��}����B��T� ���ps����I��/e:Z���o(�5�!΋Y����� �(Y��f�w��_Sv��Oɱ�\s�Qe���l\�EG��Q����;K��^�4�?�3�l=��l����в�}I��c-1L���!2v�M[D Y}.䵏�/�!�婇�� � qi5A�&R�k����y�BM;�5��a|�J��=zpf�cB�mx.5�<���TM��C���zy=�H�ze=��!�{�	�!����$g\B4��}M�NK��n����>`���+�(?kH�GϮSٺ!�ʟU�����s�cA/�0SCE�>:�� ͪd�@�u����n��jPx��.6P��u�]�,JP[I�c�@�y��/^�L���]pN�N2x�{m	<���م=�')b�M�F	q�t�k��'`C���W;o?�A�r���Վ9sQ�^	-2)NiQlGG�}�DW���$!ѕ���h�����y^-�1�
��+���T����@qt�%���
�/��l�Lo�B�P������O��ެW���lN���=���a#W;���K^�K�����f�VP7�#ϴ��%�2^'�3L	�?���|`ƚfWvD�Z�s���;.�����vP�5d�yURz|>~���v��w���Q�c�����02m����'%.W+�%�+>,=/�5d�M#����v��}&�����ёCK��;�U��*.Ww�#	��� �ތ�ץ@w}�]?_L2�Y.G�U���j��~�����&g~/o�[���������;��^��_�9�{�a $���mm� B=��;�r�s�"e��d��m�\�F�%��M3��=ʿ�E��j�L˔��5|4_������?�9ٳ�߫�u�^Ҫ9��P�B�ERF�F�Εq����:l�D��O#���+c�N�9�epj��ߓ�jF��l�N�{����5�������Af�%�|v����r����͘,�K3���@�90	���Ѭ��M�o�"`�V��۝���.����*����� �pPJ�e$�X�sk��t-ħ�O�Cv^��]!i��Efoּ�dD�J�(��w\�=�R{���q�SȬ�M���J*@�{�5��� ~� ��ؤu�a���$��>gֶ��'svf�gU�,�f���Y$fLrw
�0��f��[t��Tmu��$��A���:\�
\�K43�@�C�	9K��(�x~1B՚���O��n�^���c���Fj>�%>R�)�>�ȓVm�fS*z����o�p��o�,5��V�p�̉�&>�ȼx0�Ĩ�D�6�17n/�f�=��o�D�M3����� ���w�ZV� g���\΅Dͷ� �T��w캟���KS���c�5Dg� �nzw�� ��::�Ζ�׻r|&��HqI8� Q�EK�z��k�=A�����E{�e�+� ���W��L�
��655�}Q��j���C�����Q��=�O�/k{��cAULl�Yq��w.E��uɤB�����ܔ���!R<�l�>M��o�� ��b�K��5#�f#��ѝa��5h�P��F@�]<����Rh{l��"��v�oZ��&������r��u�h�.�h{��7�+����4� #�3�b-z�nח�R����u�9˩%$�7:��� �F�G�����X�G���,���'����w�J��cj��4���*K��@�`1�(�7������.�уmr{���g�n��|d��h>0�m���|vX�u�i�N�(k���M��J��p�Y�yy;���WH�Z��k˾����V7?��5B�O�\ȓ+M�>�=� ���
��F������_B��IM��z<g��������eOM
�K��(46�&:�����"�p�/�H��zt�1㣿�`d<�b(L����M&l��iM݋�!ڰc�}�dc5��`RgCm/E���:]Tti�ku[�T+����<�))<1o p�I?���֌��ڼ��b�X�ޝ����u�64'��[-�Zc�M�����2��T��Fh��ȭ���g��	2�� ���UmH�>��g�r��V,��}q�P�|U:X�W��ߺ��x���;_o�c�J�X�������!#�	�%&b4�q��f��Hxwni��l�@3�����1��u���5�O�}ҳ�%/�.�Y��s�g�8��A�~�54_�yњ$�t��Q��g�g:����N_R��O���É�%jA��,%����ƕ��n�ӭ�����I�ڟZY�^/u�-�/v�{�U�ǢʷR/���b��r�k�L��Wʑ�W�,4w�K��)/��DS4*��o�
��R�)�L�@w�ٰ5����Rϵ�8��Rj�rk���,J\��an?BW���9f��p��O���`!����2�T)���w�ۨ�2�&>֫v�*�����s6N�ƻ����ça�ا��vϔ:��J`��y�z�r��qs	z�c˭�q������E�.��c$�_���
����s�şv�|��i�v�5�N�����9�l��j4?�K�
��yk]�ΖIkv3:<1SuW�?���jI�|��o�_af,��61�u8�|hU&�
�(MFWM����<B��d�AT���?����� (wD�u��^u��k(,!��)�RLd �K�v%.G��g��N�êґ�g��k"�&/�t A��%J�E�č%���<��`(���]F˱�o��X�\?� ��p�����������jj�g{�j7��]�S*�go�;�5���}�g�_ao��`KUxM��.Y��>��́�a:����^���ͷ��h-�tlxQu����H�fC*�l��hN.7��bA!�����g�R�w���tg���ϧI
7�K�����n�`~1�'2M��s��S�_��ґ���bf�<-����T�%�$u<�Wp<��ۙ�Z�H�ʎ�H��:/��Ֆ��ؔ�"mJ�˹)1W����$'�'�A�� ��.���h�X��2r%p�܄��pa�G1�Ι�,aቿ���<�p��G�H|��
��̇�(�����w����Or\�	Fd`ˉ�n�6t�X߄p]�	�u���<h%3?���3�+���m>���ؚ���_F���W~y�[m�;����^r%��)�_����-��Z|���;���^v�?��b����9��<�j\��+�&5>_߉���d�Ѹ�e���n�¿t!ke2Sh�{)�t@'�|P,9��U���o�,��?Mo�Й��P3D�n>��:�8�ڿ.靠����)O'�Ie�z�3�mV�z$V"7!���ݏ�xW�=�?6�@bb�^)�s��W�L����{�#=��҅UV���G��\�1��j,I�j�ך�#��6�S`��`O�jQ�"fG�m��N|��+/W�l������-��j5�d���N�{:�Su޺-��@�S!k濒W���Y~t.mFi6����<���4b�+����6j�/u���S �n6.�1��W�f sP��tR���*AYĔw�,�bq�����&?`{��"8�[I����l�)e��OK���6�D�B���cC9�9����^�01�q<I��M�/���������=�\�����q��9�Yw�B�+	:6�͊�0.tbZ�Mdڱ����3���S��iW���SF��b��7T�!O�z��\�B�!0�vQBo�e�1.&&[�nNz!�$(��T��-y��]�D�-�\���X����j�i4q���ؙ�v�4��1�))�[)6�T�q�OO6ᱏl��j1>�3�Xބ@L�`�VP��p_m�C�����ݥ�)�\�z�澚�)�)0R8�1Q��������<���Y~oSF��2��x���E^��M��T����o��P����.�:=O�/֔�n�HqL�A����b��^�'I����st�+����c3��>D8�����E�z8wS ���S'^���׫W�"H���n���X�9�"��[�uI�4ߨf��w�n�,s�|7ԪZҲ�GJ�sn�	�> ����	([v�H`�|���u�q�7��KWG�����5����w�Ii��%%p�\���^h���A|r\�!��)Ҽ�_���n| �]Z�Ch��X�ɛJN���Oݬ��@Ej�y	�d2���`z��3PR��/���1�{5�f�v�k�m��󖧻Y�a��9RjxYL[m����Q��gHբ��/���
�8����k3#]{�X���0��65Iw�����t���0�2*�/ػ�� Q-�sA��K�	�g�Q ��V�ڡ�=����s.�,���.;7�A��DF^3w� �%��-i��+<w�V������-�Pc��IR�C�l-���'B#�So��+Wo�I����`!ڎ�:d��^�+P��F���! ��"�3�%l�j�4��#�-��X^�y5�݂�	�2k~g�S�р���΢���>+��'7�h�9X,�f��w�������|��s5˗鿎c�V��l����;��\Mm9{U�$J�b��^���W�$]�����`�vOE���ie(k�������[�����8��+�?9�i��>�! ^Q*V3fr^�0�`�ݰ�2R͡kS��\��Iٍ�>RX���:��9�D|�fG�m���Y������׮�j)]��_�
�A�i��y�9�Ș�J�p��'��'*6�y�6���6���������2�Rg�n���y��u�:
'�����֮G���{���K��Yz�(�Е�'���T����F׾�F�P_�7���P�9DPD�`�&�?��$����cg�r;� $���s�G榠-,Z��y���J����q�H�3�ÍV��k�:d��|���j��u+^Rz�?[$�H����ک�l] ��N�7�� ��v�9>E���Cfw��̴�CVX^Ε����=^�ŏ�-CЗ��*h<�t�2�EsӱM^F���nE̍R�q��8��H�l�'b@9^Ci8	1#������k�]�*��l�=��&�t�KuU��@fxj/��H�����l�oF��|݁�Di�~`*b��|�^��M���A�x��+2q��i�h�%��I��#��(|>��r�w�:)l��� yh=�:��ʻ�ϕ6��K�tÐ"x������wT^a�=��9��щ�.moO�3lR:�� ]�t��S.RY�Gh�lڏ�=#�#E���.��*��/J(�R#<>��?��/@�E1��ѽ����ƃ��m��2��T�w�	0Bx��i�t��u��d[]tN����K<*Am��ǻ���������eM����sL.��Q�$M�L!�� �֬!�\���i�K�U���:}=�_a��R�5�U#Z����֑sb�W땐��B+k[��=���>���E¿����)j�����p�0���bid�7;Y҅���6�w�}B�B�ߌ{�]@�%$\$��V��-�,bf����ޚ���-��`#|7͂ �����]�3�N��>��5q����HR�B��q�0�ש�5�l�J�9�Lo�E~��bD^�)��Uo�G�`*7#~��>G{�r�0�7R�K�m�QI����U�_��F�ڼ1T�+j%�ł8��x\�E����B�[�~k�,�E7-"���?S
d��9���a����ԬM�%"@��0�c��y�@-A�l������òj.!6HOm�p��$��*A_�sS������G|�y+�ؤ�j��i����>��7���*���sH����m�˲yg�Ml7�cm"@��/���d���j��Џ��A�p�iZZ���E_�/�<sW�0`�bt��*VT��k8:�$�<��z�B��z����w���L��v�y�u�����k��3�@�y�/��H�*+���#P_��U%j�0F\qR�/e�T9�ю�� �w#��Y�r�3�<�e��{
(�p�름a;�Ʒ<;�z,�+���K����H�:I��`�ç�y�6��~���bֆ�Œ�GR�'m�҉��GFw�����w��y&ߢm��W������ЮN��ka�Sy��j�x����9��={��tc���6�9.��Z�����u� R���(9�5���u�b8�^��R�O^_a��E��:�\\7sk򾘋�v��%�ո-���B���Ag���U��`���$�i:�
��_jP��S�߲<�@$H�����-�c���!����_t��(��nb�*3��l�8#P�n���~��weÏ�� ���,�%/��-��{43�ɚ�	Wv��h�x���ːE�����F$�>#�q�
�-1�S��i���г}	�ⳝ�+���5�x�XI(���?�c�wa���G�Ԝ����ѿ�&2��#�P�x�R�JR����r^�_���+[��k�5^'uu�R<o�u��Ogܛ�{����2�9�|��U�,�5�_��zՏ��#��6>A2���N��yi@���p�=�N�B}��̮I�u�����W;�UYH��ЎENg��bݮ�۹'��L��|�Yo�4��{퍪4j��
DQ��V*��o����m�=��. х� rDw��9�<����\N�P�rKy͓�����P���ܬ�D>��	�
/	=�t�4�+*�*�e7M���y�zKR�K�~E5�=ӵ`�Z�L��I\P�i�#��iT���e\�wxkkU����#>n^��+4]�ͬgÏ`U �	�'y[�D�e�S�U��w�>ed�V�'7���y}�	ޤ�u~�܈��$��S�c����6�Dr���!���TXW0�iaƕ-�$D	Q�����Eq�|��m!�q����=���@aK������c���AHT��� �uwa�S���'
������ޒ���mc8Ryf���~#6�sAG� ��;fh���f�9�^�$���Y*2�	�4��dZ�
]��!�VF	�NW����v��u�x�m�/��9��i.�ڈ|0�/8�<.�Ji�s����y_�{9�G[btW7o�$�,��=&ka��l}�rҚ�0
M�/�yQi�0����;4<�g{�8����Z/r����؇�/)%��Y�p;�E�I�����	aݝз ��H$>AZ �^v�/�m��!\��Snp���£�j��R��@�r|v�;ͩ����U�}'�(X���(m΁y�i��㚻��t��� �p�|V��m'��G��Z6R#$���@�$%��\�ȧ��d��L#����ߧr�T@AsԒt�h!��:}�Ob$z�����5�$=�s!��Իm����[[QY�kQ�����USa��}�X�|2h�G�c���R�Oda��+b���< �ޘ�0����*h�]ɪ!��\�m���!�t8��$(�J�5�^�Y�o�-()@�q�����=� W�X���C2����kU�%TN}��N�k��� ���x�L\��䄒j�����	C�����y��e�U���'��N���D����}b��_�n�t����.�d~�$��I}�c�3�s�W]�8�@H���i��@�V0m��Xr�“��j����X�4�#���Lj�a �B�i�^xK�+��hO-�t�cNr69��P�8#\�屶�l� �'�b=a+�N8q�EC�3�_*���N�ؽ8L�a���a�'������-��7Gۆ{]��� ǐ�Hoq�T�'�"�Zs @�ט�y~�%;vz�1��A&L�8)`��Ҡ��\�
��$%]{�0�b�o���ۧ���x�đ��!�f�u����¡|�I��oХ"�ږ�^ސ�o������kn��������D��U��Sg�y����+_6�g}X,P��f޿����F������h1���%@Rku��Dy�'��|���(�,�Q��<,�z��p�'=%v�L���G�7�nfC�����l�v������
l�|�����}�F�r��tʑ�g�	%�~/��"?�YA{�`K �X�k,A=�4���+'��H�3~@�������&u�˅�n��nȜ���a�e~?:�]�D�M`=�0��h���ԣ�[�2���w�#C#[m6I:�ɪ�����ͫ��P��-��I��P�,�g�N#N��R��(~�XlxV64EB    8b3c    17d0�C�w� z�1��:L*�U��h��[,�EZ*�pa�3����R'`��2`�,�!���3�cXLA?����('F
�[�&P�ѶlD)��7E��kˁX������:��w�u��-� M�Pg�{%�c�ld"�[�s] w;�����1-F��i�68���HʀBu�j���lw!�.��HD=�o�[��Q�%�&Q<R��咝�Gtx�8�<��Z_zϻ#��soC���r�X+u���2;�h;L�����������o���g��KȐG��$p���Tn"���&"$��YR�b��Q3R�e�t��X_|��>gt���d�h\bч�:�'�"_�Gba�"��pX��N�B�b�i�µý��-�`�P�Rc�lW��t���	�4���}b��rIl-��-}����Zu��[4��4���\%�0�Ё�`�NJ"���[�ӂ�mt
�EE�.z�m�Ʈ�_pn�!1��'��D�v��j�'�wuW5��W������l%Wmn@뎢( ž�ދ%��ps��Ol��4� �Hǫ'/��}�|m u�j�or 6(���2��06�qH��#f�Y3�����d�9�ɝ��kS-�� ���?[W�w�!�²,�A�XE���\g�Gd�9"����d� �i'����W,kh���������K��~	�ML_����T����>��Vc(XFTL'}|M�����}�;�Иߌ��:r�1�z-n�g�6��h��%���8�3��AV��
<J5sB.=��sI���������� ��lxr�s��}T$��kk���y����QS~�/�z��
�d�<D[�9G����3�t�rϗ �(�Y����D�*?�R�5~�v&N�.7�m�N�䰞N@.�Q���|��=��3j�pO�����	s�ë~�3�,���%]���١�J�m����l�Ч�Q��V�{�C��K�U���P��c���e7wY�~�r�c�`!m��i������g���>���Z����x��#�4��W5��ۢ}��Kd�B�z*�w�
�Cx$�x$�I�� ��xA�tO��z��*�!nf�o���*��=�����Mj�A籊4L�,$����ڂ� �^��_x�5+!�a> i`0��}qE��.>�9e�At}��/�7�]d��%����X1dG�٦���K�۱>;��Ϧ�(����5�\"��F|��_U�)y��hF蟬&�ﾺ�a<�*��n5�n�(]}!Lz��eRWY�����c��uI�JD�Ng��m�b��(	M4��(ו�f|�"�Z�n�W�M�$J����˱E'e�FF�~6��y�ִ�� M��߁hj�Ia���f��N�j0S}e�����g|��+����#Z��kJ���fGli ��/.�?����yؤ�R��O�����2��=|T�f��d�����i�'fC�mH���q�"�����;w�3�-���Qȩiiۘ_ ��L<����:TE���lI�!r뤔��jdI���U�ƕ�1�dw.������[N�����n`ۘ�u���S��J P%���&?[�e��RwJ��gR\[$kS�_
-j~�V��7��]�r[)��1��ʒ� ��g�{�.mrkq�w�q�6��K��alq��7��f�ݽx�3�z25��7�Y���k��}��h�ycj�A3��  � ��DM�-���ҕe���H ��¯�9��|X룸�8L���S�$����y)iG(���~<6st�]���t�z%��
c���J�O�A���踋5x�s����\�n�C�/�?At���[�N[�	]v�n�!,�y5\MH�SR�[Jۿ2)��1<e�䔸o�9�H&&fE̚��u{16l)ܕP�0L >чb�]n #������"��-�oL� ��p��zس����8��g��ʎn�8 9|��K�ċZ��d���Cjn�=3V?���&z/���l;`�xQp�u���8�Ī7�E�WGK��n�C��8*\�W��̵D��{ٜ�^%�_�@����~�2�8��K��ŉ*U�ʝ��n��*Ao�'7��p?:"�a{�rp5�7�-���ү�Fp|�l�"�C��Ɏ���M\�z9op�^=1���\3,��t�Sx�2#	��)	���WВ�nǽ��BnD�e6$��,��h���h�XLV��kЈ<�V�a���>o�%6y|���\,G�1\Z���5�=��-���ٗe�{ Xnb���!'��~?R�,�ID��:�9K�����\%5}`��Y/�� a���Ɩ^����Dm��
�β�����*�>JM���8ȁ*Ӂ��b�����Y�8 T<I�ƌ�,ޞ�>��p��AI��|��)� �Π<hW$/��$�:k��v�4����f�0��2A����|���P=#��!��O?�+� �Z�Oj�L�"�k����_kpwz�X 9>κ��j���I� �u�ӸRÊ#����.֩y~(��~׭�a�/Y6P���,"?in�����-��sS����ϑ��?:)�+��>�+Þ��`��Ut��`m�<�[h/؛��a��,^�6��$oK#R�9�n6��P��kV��Cr������
���G{,��wVd�IP�u#�CY����Z?�G>�:�pX����� �����H�]N�OGSp��×��D�U7]��<3`��ۼF��F��`��[;&D�r�\o��S�{7�و��l�F���/���MN���␔~��C�~������ަ��{�Z�_!��[��3U�Q4]��-�:����ݱP�6vC��@��坦�V�T��E	�#0��A:&�kDj�_�I_<��Q��"Gy�&�V*��N�z�tЧ��*^��z�����ӊp��w���Ë� m�;�m��1����k���pA\zU�=������'F�����j-%�PH�����^7�Z �������#fCu��AKؾ�����ف�w �Vc��S�^���KS�^�*��c�!�WӚ�^�Po$�|���ә�:����bGn�0O�M�#U���SN0l%y2��[��a�
��_޾�؈��\O��t.q�(�}[�U8H��Ɖ4V�����=��f۵/�Cѫgx�<��S�%��?�M����h���(g�
�+��)K��l扨y�P��T��bb���Y6?PԬ�,��)���-��������m'�یY����З�G��6wA.^e���Wnҡ<������a!֞(C�҅6�V�OXӛ�}P߭:;�)�*��v�P�E$���a�<HMW����Is�D0S˩r�p_r��(�&�l�=!!���-�;���T���c�+�'���mF��h5'8�;�6�a�;u�}��nd����~+�t�|d�ޞ��2� ��R��揣�µ��
�ftD(�+�8�,�����:��d	���2�ҧO4�3����$�Cf-�*0E�TÑ��u�y��\�B-�n�k� 27b�A�Rud̷E��|6O�^�e͔����8�0/*&���tK��Z'�g��"6���4�lC�e^���� n�X���	�+����%� ,�|{URZ�'���&��z�Q�T�Үk���=���_$`J�v��Y"Ly���s��>�e�s�4�;A|����Z�%��V׆ig��g�njO���;y���TxXq��82���>�3��%�JfGل��ݾ�����f{��7e����A��z[�(y҈��	����[b�/&���Tlz��40�Oš̩��B��12"K|�o���׺�\��p���Å������6�~rzS�*fPJ�Y��51}�ϑ>qa��r�bo��YiDE)y��KD{Q�kSL4z�Y��,Y�,ѻ���?��U�R^1.a+�q����:�<�ᩓ|�t���G�h���=�e�	�W��2�<��9��mo2�J�Qk!�W�
&��$���6f)����@0
��yF� h��S9O�KEMS�"�2�'�����@1�� �zca1��z��K��]ˁ�S�/�����L�����C�E/��I�~x6�����)����K�V��nz=X�m�l2��q�&�Ύ�Cz!��sB�N(�^�%\(6�H%��7R���hx��~2�s���.l$�Ex�"��}�m~꯾t���}3��(���;��C���ٜ4��I��n��NHV2%>U�H1���Z1����
����(5z$F|U�ѿH;ztAEFvhY_���E�OBh��7���4T[� \+j���ڥ�33
wFD��'�\�D����M���R�p�񧳀Iaƹm�[Q;%J�gTF����ك�����"�>i�C���b$p��\��z�[��F�e�#��qFĻ�~	+	X,QL���s.��
�5i٫���u��E1�`�f��*������-xS�Yχ�#35�g���z��f�C\q,�^B�9}�$܄4�e��$��[�o���˙t��������X�� ��Ku�����Z�),�像@�Kג-�%h`�H(s�K�~RՓ_��?W���U���H0��ʟ���I�OM�B�w<�3mm̮��˓z'A^���m���FQv���[��~�be����a8G��$"�"�5�_���%�.T
ܴ�����S[���v�C�e��X���e[�;�A��+̝�m���}d$P�D��鳿a��"<9�.X�bD��^���x��0����esP�iZ�ʒҌ�]4�GȳZ��2�e��/ڕK��A8��a!)�X-e>��^~�:���A�
�:��i�9"�H{�|���ĀZ�#�d��B���j��ţtqE��j��1��C/7zK���PN[�+D	=�u�3=�,o��EJ��e6���8���Q5(V���$��ۺ4�q�n��|d�'��:X�L���J �rJ��&&�H3q~��c
_R\�ݙ
�~X/�J��w�;��S��Ѝ"�n5�o�Qi"��X�R;�eh�T-d���$�/�k{�&��S��.��4W��큾U.xlE�w=��b�>o��6�y���c	�&4� d\CP�N�R��Z�D{�X�L�xX�����?l�����T���l���?�˳n7NC�6��D��)��;�+Az�D���{�,�}x��͹�S���;�)���['K�Y�}^�Sr�v�U��C��8H�1�1��	f��Hr�)�rω"`G]U@���F��H��;J����B�DbE��)�FF��no�.�eHI�k�guO2f8	���uY��+��:KR��tn2>��&��PX��8�E����@8=񔀕q�����P������_���y�S��y�S^gت��=�T+���a���?71�}m��4� j@�e�B�
�pTm�����f^�y�=$����T� ��^�~ܝ���4I�>�����RX�7.��ÂV�'����49� CqVXv������h�IN���L~��e�l�m���H9�0��Z&�]�t�v��}���w��?<��u_<�r��Έ6m�Ͳ��?��|SA2ޝHF��z?��m����-C7�+�hR`�Z�ͤ�$����a�A
��>d,ɇ֏3�׃�@9�V�}B��16�KE%�3�)##wec�|�h�z	!�W�˶�%�d����7�dq}��S/���A	�B�	�V����O_n����G��/�l<�&��b��,�\����S����׀Jrw�C�c:z�,�dKi uSUb�ukV�5Dd�m]�������E|Q4Dz�y��rG�mh����.3Drlz%u;:�������c�y�V��mo,qS`��f]�p�WO��p�Y��`���F1o�u[�N��kX��!U
�\�%7�i�`��+3�A���X���q��E}��*$T�����a����*�F�2��;;���Tt)F�
E�;��Z؊�Ri�v+N�O�$rT�,��n#�u^�9u͏t''�w�}�ֵ�uf謣C/