XlxV64EB    1825     990�+~E�@��l�B�bt ԓ�S�-��7<	_�_�E+hw�弡).x��t]�Os�@=��<�f��Z3��B�+��U��t#��ŭ�*��\L"�6n<��Rf	Z�B������u����V��,�a���ru#U4��c�� �<�m��н�WB����؋�]�{{�У���xD�=P������[W|�ۨυ���yyD�A�`�.��"iN��æ�S  �n�wPh���0��wr\�}�R9M�j>�ǚ�P(����Msy[��D����5$�]���A���7�u����@+<��%m��pSB���}�Ñ3�Z��
��#�9���?*v�����5���X�6#��6�\���L�-�"&L�̲���&���
^��F�� Y�E4өS��,&K�(��A{����j)�Ui��p��XҒ '��%�����]�Oedoqr�� �|�n,\����&����[�2�~����� a"e�c�*��L�X�����~  S�q������z���FAf�XwX-�fa��@$�y0��\��|�m�� yn�ʣ<X��0�R��H���?4E��8����ꟇC��t�㽸�������V�n�a�ﰠ����^��á���b�
S��@�K��v��ݲ��K��s��	@-��5}y��R8�I��M�Y�ʎn� P.��k���R4Jrbb�Y�L��E�.k��h;1��T��b Vb����OzT�v�ڤ?/D�C@6i����1R; ��̯ڢ����&�ׯ�b#8�#�'ֿ�^��"}��h��2�x����}���bUm��rW���c�[`.ή�
�C ��t(�b��fG�h��?����fV��;k�W�p6��_(`@��H�)ѯ�����������<k�ߠl��op�x(���6ގ)�C�X�U�-*xa:p�x��l���o/�M:�g�|M@����"1���yP�V)?;�A�_�5M��-���
[�MMIV������N��
��E�ɅW�"�o��j��Vz8dL���۲�%��7
V!�ѭ�%��A2jlqΏ��|��������H�D���H�`�r���ۓ�H.W��+��@�d%��$�aJ�|�G��V�	������&r�A�G��X�l������y��7U�:3�ڳ���w������$�e)�$�f-:Ѝ(��Ck�G�I���^��IJ�k~c%�}�Ԍ��N�q�y�%\����:
 ��!a��GWJ r�#{�)h��;>�qB��r]{�&�6M�_�*GL���G�O��}�&�"/�$q��Y�NI�+����M��0�>���<��e=�a"^�31,w��܈��ԻX��q��^V�A���>N�=zg:
�
���Qs��^�"\>C-<G��/��toqI�G5�G���bx�'����B�=��@\)U�l�$�����Y���QZ�'�*F��is�ŶJ	B��A�=9r��s�o�/���_�R#^��I����Ԣ�4��)r��8t��<D��O�'D.H��B�+�z��$Ɋ�v�&��(�r���ֹjbL�%.�Z�Y�)�$�W�Y�YP�/�������4���f�vF�j������v���M�Ի���>s������y����t ���"��@J�%7=U�F��ƍծ ���aU����j��WXh��������Ԑ�����N1���*��.u� ]à�
*-���-�^:�����U�)g�X��Y!Z��x��k��ԱU�B0��>�<�R��q��0����{�����ܺ�m����{����B��O����&A�.�2�9��C�q!(,	{�w�Tj����+*	h��*g�	po�9���(��� ����F�GeT'^�uC�"�X���А�Q��b)GJP��%��K��iE�c㤂�Fe�����*!�?w+��jĉ��ޕ8��Ç�j�������s�ct5 <��P_2�iɁ3嫡���F��#lQew���iG���Skf����g�w��j-���c0��o��CR�]^�A�F�HN�߯ks��K��%���OA|�f�7�/�ۨ\:���<@��'��!H|�vVU�B��������5d�&~�����?��ң66�J�����i��.8��祈i:������{�	G���:if���m`8@�]^��Q:��L�����ڙߏ �Xc;V�U6�]�d�"T�ꊞ<��W�:�Q�W5e	o7��=7�N����&�9k��(-!����ʹ�%\�T�С��d7����:Y5A@�&$�H��Ȅʶx&�	�ȫ�3�I�b�"��s+�Q�M؏���A���Vx�"���L�!�����Y���#X��L�%���?��C$��Ҏ�a���A,�H�t�j�;ʫ