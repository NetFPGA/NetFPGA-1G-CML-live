XlxV64EB    4336    10c0�D��	���X�L|�7Q�q��9jR�!�x�� �3y�d�5oQO�\�w�4���ʍ&�WF��"�*X�*�E���{�s9ƫt:{�h���(B��L�X�h�n�����|����C&��O��򹸇h�Ĉ��M�Y~⌊���j�*�UŚQ�Ц�
�Cr@/�s����d��ǻi��-at���7sd��Ƃo�;D��3��c�>$el�|>�f��bV�諞Ϡ�5S#�%bz>�c	ʷ���I:����X�t��rzy�Sq�$Y�s����L�/EG�Rg��BH[x�]�����kB���0<V3֒l�����-����b\sv���9�ⴅ��Zv�����{E:]��є� �À/�ylP	����FGŊkهm�@IE1�Gzp'��[l�j�*�(�8at:~R����O��㊱���*Z�|�� Zx� ��4�t����D�&￰6����R��+���� B.�#�£�|�t@=��;�[�'��?�6ڱ 5����$RGM���˳� �T~��,� �C֎e�R�i�id��C�!f�19�  /�ͤ��sv�e#���K�>�@�0����4J=�Pv��-*�.�#>??���!�ʉ��	�r���xt!S��ɩ��`��OT�p�	���-��mn1�s���}�<d�-7�U�hq�M��K��L�:��:]Κ�2�X�哟 ��\���f��E���خ��|�h��i	|��OV���l���D���V�6� J�tvf�Ү��C���S�����=h�H6�������<��7T6l#6�2Ǯ+��%!I�
��p��]� NT��6,�7cr��k���㒎�8�	$ڗ����59��/z��;H��h���vŔ�)�H��b88�B�]}��ڮz�?���=G��T *[a��uO�[Ω��Kud\�ʉ�c�[�a��Uw��+�>�ʾ��T�bc>!����e�6� �I�D�U����,"+��{M9x�>�G�p�	�[�^V��2@m)��:��Ko�#�a�Z$�d��b�N6�W���8`:��a��>Y�$v5�M�����帊����bE��^���!�ԁ
Nt��+k � ��3��4ϜY�Wɣ<����� ���F �1|nE����`2�Bg}4s��14f0@m�1��x��1"�ky��>����lFs���.�
D��}"\��K��8�ӟ��b�Z�N�[R��3��c�o������zf�wj�_�<|
�J���)��?O�+������SV��\A%ƞB�h����gu���Q#�(�⧻�k��W�ٓ+���'�"��F�jw�����J�_k̥��x�ֿ��L�EE�� �����y��t�S�J��,i�	@Bex9�8>4�x��,0�ⴜ�3?��8�
{(]�~�5��G�K]7yԶX�ɏ���#����<�H\z���d�uM�U}:�� �U瞎��܀Ҵ�i;�m&:�/�<5�M�A(�IwK_��a�''PT�h^���&���J���ˣ�9��,	߇�pK����1A:�]�"��wH/t���V(��6|���7�ĪL�I��n=C�����]�k�g�v��M� J��:��-]k�E�<�#ב��boQ�>i r�b��+'�l$�Q��頙�o��A&�kq�3��ŉ�5TY�ڜ��Ⳋ�Il*3����8�>�vd�_�{��u(Jl��D�B���q�c21�$ݕIw>��;�=���j���	�|���9$�1�	���X\�Roe�ACΏ��Ga,Pb��$r����E�����f�JA񿶎�����@]�����������jm��l�]~x��%�WM"�f�4#��,b�vf@M?���G3y@����G�t�� k���}�9�g#E�S��:mةN~�?���z��U��S��x�sp@�#��]��!̻^�`l�΅d̹~>�o�q�{��>��9W:΢sz�ð�h-ڜ���F<��I�� 2���D�I�\C+�|�Fy���]��c�O�<:����c\JH��9!���4p
�S\T�O��e,S&����>�/��첝�=+�/��9��6R��DϚ"@0��7OY���=8����q}��� 9�/_
�{��%E���/'E]$���ê�>��E��<� �����QUw��
ft��Tj8�:����ʸř���H����n�|��dL�D�r����y�j���ڍ,�稍�;�x�ꮃ�q�KBE�옩�y��m��ף��7V�t;�A���̼����=��j��H)	�R�ZXS9U"�]�Pp�;�/̥�ʠ������L�O�H�ǰP(%W⮿�M6�����~S�����~�F��%@.�BN�Vj���	-?����te?�#4�R�[%��tP~ؙ�$f�}���]�U��ԯ3� ���kQJi$�Q涫�����]m�q ��޷��I��
Q�b��a�=�/Τ;���)��P�I���`s���E��|'�D`���^C�(�/c8��2���x��HI�'�9a��#�#���R���R��#��P/��5T�m����STˮ�<Y��p����̂z8V�v��#bS@Bd�CD�{�� ~H�lW/�%����?�qp���=�bHEˉgd��\
3���#%Y�N��`��U�	�/������
�	`}�T����-������Q��Hg"յ��wK�`Xd[Y*��3�Ԓ��
��?�G)V1���4'�AO%����x��5/!.�܍dO����Ս��C�Q|���T��!pu��SЏ�������ۏ��j�?B��fd+zB���C���!lW.���ܫ�6�z懤���a+Q�����Y� �ܰ�=�p�v<�
Qt�^�R�r 1�\�����}�	Ε���¼Y�����m�qv��\�j��}�t���X��݊造���x�_�Lq�9)��JB�\]'�I���6ֈ��_��#�_5۲ѽ1S� ��{?�0d��Իku�@��(��@�j�-�Z�m��p��	�WtB��r��� �\��J��I�hP�=~��i!�)��ŉɸ�A3���`��G(���DH[S���rA"����v���9��GH�+�7���ܾr��wҖ$��6�~�2����AHk�N�U�;�5��ŉ���$%��}雵��������Wl%�ԅ��J�įE�8�[���'t�_��_���;�#�&�]�E�Ș�d��` �S釴2�DT�p��*��ܕ_�7�G���,������̵�.�f?ѡ$�^�B���F����F����^VB���ឭg��Է��@z�Zmʞ�%W��������$�(��i�}����z�)�a.<?S�z�KiY=�
#]�%vS?�����=X��	�j��[���ȏIb��{�����.#@����ҊK� �>쭖��T̍s��P�B[S�TԮ�GEg��ɗ�����,`?����a����������ߐ��+��4�F�GSn#�B��/f��v�j،�\=�S�ު�w����D�0j?��^�!V�#��wJW257]���?�Z��}1.�{qiB��i�?��U��<8�.)証�c��<�1���h*��T>�h�R��97�X���ΒI'�)�Fsn�ɩ���І"KF�0���0���exO���PJ�C�K5���KY����8A��(�X]����y v�]�<���g����>�Y��[E��~��a����~�]p�΂�gxv "6Փ�-S�_o����� � !Nb�X������Ot��85��+}lT;�6��.���II;��G����1�x����o�Q�r��t�vvM:�ګ�1��`HjȻ�60z ��������5����<�U=~��9gV�x�C�����+	�����
������$�7RmÜ�$���18�����$�c�g��LB~��#o�V��}�^�Ol �̬~�2�=#z�b�=c/7�y�kҽ\����^�֎��n_�����T��+7E'L�y�q���m�*<�!�7��{*���f3�#��߳�hpz}4��w��w�h�ƢA-��ik�z7=�p�Zט���Ro^L��ԾoP�*֊y���x���4>c�F�ѓ��* ���8I{-M���nC��9p=�V�Y���x�-_LIʱ;����q�2B�D�h�=5�`�Y�