XlxV64EB    4876    1400��(���C˗�ř�PbY:�&L��dqg�:�G�*���x����7o'�}�j�Q����6i��"�. �f��38��g�����i*3�����1�vE�	M�4��.^T�4��G���?asamIJ���g�e�����"1�w�5�=щ1�Ѿ:�$�=�,}Th�,s���d�C����[���D4b���U�׶WI��J�M�~p��0�_Pz �$E��
10� �V�A��,{R%��%YQ�� ����iV,�P$5��!���=��`C2����4?��_��k��/���v��v��9���.��YVΧ`�-]�~i�D�n ���-0���aV�@��}hT�e����hU������r�����m�@��u�����G�| �x���fD��\�z{7��M��}�)om;�Fd�o_T��y<��,��Z��O���@�n����*2'�KgC�<�}�+\3Ƣ=i*���>����`���=��<[�pG����
�e���#��a�L�[�5#���E�&������* P�OQ�0����,�,��fP������}F�L���k���^V�*8��ތϷ|TO4/6s�h�ߡm
(�L��"�e�x�'"��^�0��E�F���1R���S�q�m�R�����c�|U�;-ZD5w^�fEx�VJ@�Aް�6���:<Զ�;b
�}2� �UXV�oTW����� �@�\��x�>���)�EgB����L�0���x����d�Ô�)��=U����k�!n�sU,��i`�{y֕Y��_���;��J��ohEp��t��^#�k��I���=�[�L�|��$g�X�B1
����˿K�A����5I��Z)�7�Q�CK��@���b�J�G�[*��g6����o�AG�����h�k�;���s�DG܃��A�LpƱ'�9Yp��}{}�e�Io��ЙC�\D-���"�[/��ac���m~ƨ�5�H��1,��b�H�Ϻ�B���c�A��NLg0��-h��M�6󆊧OϽR\H�e&'Z��c��`�i��1d�� \��-��tK40�.PΤ.n�����2���n �[^jO��1izyc.ПX_�D���J|���%�����י�GU*V^�ϋ�(�y��Ba�e6�p*���8c�|֯��(i$��n�|0.�m�{�+P�J��:��+��U����Hg2 �|�bW Nm�k���JV�\E���
��bn�h��9zu
�N��l �B�tqx����9#�b��d4
h��7�>?Yŀ������5����i4�wc�`�Q���T�hz�G�59*�ײ	NT���#�%�SL,c@��ፔ�ZV�z7�[s�����R6�#��A)Z�����E��ٴ�O Wg�-("�����{sC�y7�VbqSa�(���괂�����O߄�uX�{A��+DH� �F���c!CT(�Q�?b�SXt̪|cF	2Y�Fo�D�ǐ����H��&\�zI���Vg_H�u�ׅ����ޕ:�0�{hh��#�Yx�ı��-���ѭ#����ۘ����Z5b�t�������a3&��RL=Xlt���\諭 -Ӛ뷟T{�N��!�л��2�-4�b���������yQ-6)�eL�=��<t��k��Q����N��^D?�Iq�6�:Օ��g,�㵩���r� V#t`���Ŏ:����H~ g�]�z|��\�cA$-�Ť(km�C`�O<����M)R���^�'�ut��¬�v޳ZX~��Fq�e��*tӖ>��KZ܇� �t���I�M�1o��噓���~cq�7����]&�!��G�q��t�\$�f�Y�2o��V�4�Sy�du�N�@C;3�N�)�?Dj�e<.|�8��Ώ����e�!υ�����+�2�.��/����#��^�XMc��r}`1�T5���-d�NgW�\9���߱��y�H$�)	M������J폂�u��_}~[ѵ�Mn��mB;^>Jܺ�ᨽk�ǝ��(���v�(�+Ĝ���Z)����e�K�����S��N=D����������"��FC&��ݔ�t�Qs
�v昑��b�:ùX�x��(Ih�%�t܏!���:���/�:f'xaY�F��A���Y>�]�<	�1Ⱦ�s[������<�R x.k�����	��f�a������'!�t/�%`����e�� �?y�ǭ��З�ʎ�U�d�,�w�sGǪv�ֵS,���x]�2�����2E��)]SK�}�vl5l��M쌀3�x�0q�����E�4F�O��*���`�jG<Ձ�1�T����r��9��d�Z#R�W�=��=ܯ_�K��j�HUXj���ߟ)%k�HS��?w�jέ�����̀+;Q�'#\�k�ӗ"o�=)wpTA�l]4�Pcِn��J�Y�^˸f���Z�)�����W�]�>��#i���8�J�$SNꌆ*6X|�v�o�5�Dv��C�4�;!�3��=L�@�M0�i�`_f�p��.��)�����3a�&��0*D�5������'�m㰙p�����r@pǫy�v� ��^�6�I�84+L�ͤ���Q-C�]��y�39��%����;���*�����]�6<ͪ�xW
/�l�^�����mN�����Gj�R�2�� �(��u8TL�%b8�+�g��#����#1e�f遴���2Խ �P��|J�N���L�)����E],��OD�psIҌp.9�X"�t��Y��ޮ�����������!�Y[I}
���nF�,�^����6GZ5�n�@=�ٛ�`������(I4O:������5u�/��C��7-�@3��֑"1[a���7[����s��!���X�4F>�MD�&��^��k0�I8l�H����6xp��ji�q�l�e��p���SZ~\�ֵ����`�4�hKw1��f��5֡��b�A�����ëtK_�)�{%�:�م���a�U���f�>R�|��[ۊ�tE��=���ƾ���s���)d�=/�{�#=��zA&.p�i��dS�6�a�vK��:˙��"��5`P[c7 :~�C�"v���C��Z�?	$�|`X�e��>�����uZ9���������[�e���I���o)��w�$#�}�����C�p��D�P\�k��3�]�u5e*�82�AŰ`H�?��A�9�Ȕɪ���Z1+Gɉg�-3��j�<$����m�b&F�k�*
�683���I�=���U��?�����5��06P��UK<
*�tu�ha�(K���b��ݚ�����s���ݶ�2�]'�"�2��4���#Ά�F0��K���8S����.P���Xey>�����>AЖNg�=$����)ó�&���I������hL\��+f^���"76�Pm8���%�
O��v��7x�6��jx��_�8��@ �#��%A����&�
#���&�V���꾓z��qm'N����_�c�.$ؗ��_y����5�`�y,�Z ������\����s1:/���ԋ�,�*�]�w0�qz�����@/���=WD�4��JQ�R:����4)�j?TH����-w�|P	W~�;�H1 ���[wJ8�ܷM����Hy.�5�I躉�J=L�֣�H>�x��u�(�.�|�N��.\��S40�A�"H����J��,�[Yz��4�۞�Ņ@�`����,��w�){���V*�|�;�;���@Q���|w	:/&fV(�aފ�[�����^��
�BUe�Ag?���-��3*�1�_<����jvՐ���~ &a߯�A���I#��x��-S-�{�{nW���x��W�J��/}���x�h��L��=�		��c�rh@��m;?ml ���m��?4T|�M��D3J[h�Q��{��B)҆,(�trӅQ
u�~æ?�v"��Њ�Who	{�t�gLf֯��G�L4+q+�ۀ��B�hE��J�@zV �`Ë<�PF����)ʫ/�N��]J�̞x�sp��d�[�����#�@�@�`t�x�)�)([~#�,�`����W���s\6��z�|بwߙۑ��,س:GE�D�����<��h@M�Z�kU%^7��.��w~>и��(X���������dl1<�{ǖ�0���1��O�e��@���E����c���PM�W�����n|wN�����U�CÁ'-VYY��C�7?�6�1�;�$�� �P��/���̖j|��T���t<�����%�vR|�Խ�׮�/�,�]Qy�ݫ��;�y�=���K�"�8��!��kk�����">��S�b��N���xܴ�_�G�IjmUL^�F��LǤ����A���L�ڟ��M���Zo��Y��rb|���<�qܑ#/�i���]�� d	T�6�X�T�N�a�Fɉ6���F�N�,�%F0��dh�s���yW]�6�/�p����<�e@��<'�����;˦!���"Z�Ƈ�Qj�&娢O�M�+�0�1(�f�'5��l��
�BD�t�5֚Uw];�+)�I��(�b(�H��~F����nW��ė�>�G"�~�h-��6Q=��AX��;���Xߌ��A��eIc/J��7�i�_�>-y�9+��`�=�V���	#��&�} 3���cen��O�!�`s�d���Y���EPO��Xs� �y���i@���*�d�:��Dg���u
�d�����6����61�����q3���h�>�>(R���HCL��6���p��i�C�ܴ�mٝMB�J����k�Y��D�z]�p��/}����\q=�ɺ�z�5B7p��x��D���M�M��R�����f��"H��a�N��h�Y�sې�;A-z�	���wi�\�oM�;˕�ry6R�U�u�zwǇ�%<�Z�dᨕ�(��f�t5.���5�VjSF�_Er���6��_��,��˒�ۍ�D
	x��c[Q�E�<pkJ)�o�D��X�Ib�f��	x74{1�= <�Hu��hs"yޥl|��