XlxV64EB    5750    14c0fh��=8p��y�:ց�B4��͙d�x�Tu~m�W�%<��i�GԷ�=�&���ĸ�lGG�B�U5��=��}5�#O����)2�W�H�Xe�p��k�Lr�>D�}�̅�m��B�52^2����jd|��t,Yi_<��I�s8" �̞؅zz��p���N��ND��KI�t:Y�Tr15=�Xb_m}�Q������g0p0�ˣq�I܎J �g���
x��9!�}0O�(���"� _w�����#:�R��~�v$2Ȃ�xe�x%���>�Q��ׯC��pc'[��`�_��f]��{��]R�9y�(��a��[��(��[�os���5��O�."�1Udq��S:�[�LR��?�e�=&7\���,(�wyw�� ��0�%/�gɺ�P�V���Ί�*���(����4�!���q˩}.DCB�l�{�އ��UbJn.��$#�Z�a�\�$p��Ȉ�T%X�11�x��}���{���a���M[ٗ�5�A�AOFʖ��_��G��SP��>=h�F��F�w�/��}SΉ��:�i��ES��G�1�X+��=Y�ʰ���� PW؃��^�S;z���1��>2�j��bvd�m����vB[����!:������z�W�6H��ϻ�	K����#�����e;���O����g�6�(��`��o�@R��i#T���$�����\B 	�7I��Z��¦{.��d��tԬ�m� T��XHl�������!/�"�"�J����*� �z8t��dU��(�Nb�ll��e;O��F���'���d\*=��N��Q;5�h�<.��t��`��"`�/�}�AXY�<A@�+=�}�m���uǪe�_1X����9*�V5�Y�P��-w�h}�p�d����w�M���
���·�Ý�h7V�̦B�t�ƙF�z{���#��|%�H�i��ʔ!�r"�].�;�7�6�`��F�C�y���8��k��)#[��!gL4Pk�I�{Í,;��K�ʰI�+�H5)��D������r�(Ɩ�<9�����I��:�@�R��E{��
��w�+}��Rv7���>��`H"( ���T�W#�����P�$�,��Q��*�|K��+��+_7�&44�Q�p�@ʟ��e��GWALg���C���dU�Ϭ�vtD�v��&fD�K��i�n7,.�
�$J�:�,8'�^`NT���*S찿DJD	�����3�X$[�b�a����e�42�Β���t�����v
(�eW�ɕ_ct�a�wu�ՅUDU+�K&f5\�D�X�&�[z�]_��k��PL§���}ާ?*��̀e�WѮv����h��'�5�í�c����*������[0�����[�-�@����_�f)?�9��g�,xŨ��������*�E��)��k�<V�@���fuB�񫋮��z��$��!XPb�`��S�]�I}k�Nq���8�C:ƍA�����z��`�z�YZY_�`�B;��yxJUJg��CG��"j3=DT|�o�Ͽ	Zì� ��H�#g[s�R9b�nF��B!�>=/���9�f:���d������,!u���~�mܾ��RKE���3*��_�{x�v���i��ҩ�`�� V�h�n�0(2sT�������D����I�=a4��&ܥ��{��I�=��H��:���#�݊� pl�D�G#ǌ�ŲC�d��p/�e+<zw��a���^�I�`Z���Ħ�
��q��(���t���������"����=`���p`TL[��Va`"z���_�[��|�_�SXSv6+#,6ֳV̌�K�l�� Ʊ �0ڃ��X��Ҋ������#OC�M���B�o����Lm뾵[$�����f��|C�uJ1;��sv��@�S!�(�}S��8�����ӄ�A�o�c��z;�t��Q��d�ܧ���oyC����@m��x���tc�o���+��|�<\A�.^w])4 a����$�R)�j�%�_��̧!O������%�s��Ʒ�֐P���:Ε��1��ɺ��*`~8A�N�%�;3~��_=�m��z�w��~'���"��}͓Ex�<,����f�=wn�����S�~�d���-��YXD�R�¨��kj�)�Ū
��16�� >��(��q#}G��i� �7<�L�.�Нv�u���wo��
�f��{�݉3%/�V����$�]�b���+���Ͳ��rQ!_�+���;�_I����1:�lOD��I�tx07��Ƃ��� x.��c��N#�X��3`�iŘ��߀81]����>RIT�P:R ���/RպJ �ͬ8mR��b��������\��!2�J�#����6�S؛�I�8�1�#	�}e������ߣ�"�%�AE���z� �f��X�4�� �n\֖��{�o�}C΀.3�q*h�GzE�'�c�.�U�^�� T��x�	������%<��f���&h��	{�|���(ݚi�k������QB�	�!�$��r#S�f�Q������Ł���r};�,@�5��)�X6���!1W���+Ƶ�ض�D=�ӵHԡm��yXl����':5+�p.���-O #Aq!L��.�-V�3��)lމ���.�:k����0]W����m���������qR������gL��Ւ�)�ǧ%�wM-g�a�A	N��F����Q�gM�?���1���h5�"&Vy��z/ݗ�,F��.Ʌ�R��S����i�-�Ψ�*�[��U�bP��DGW�f\��Fn-I�	���U:��"�F��|L0�I+!�"����s~:Ҡ,
H�(�R�T��NJ��!qE\u%�b�^!�Jٴ��Y��vLp�drG�v�y{��0ل���y�I���H�GۄF���MG3Iw��o�w@�6Ў�W&8h:�j/~��6/o�]����p�DG#� �^y�D7��rx�-�R$ps�g�S��qu�I�#0[�g�Ƞ����`	��t25�ZJ	_v8�t�%�t��;�؊��U�$��Ԋ}D�B���������!���1!�6��^E3�\�����Ǌ���l���P��%?뚕����T�Յ��|�J�W~J���r�B�N���N��&.�h5؋ʣ���K�mP"[8�[( 
J|��b$�
�1�~4L��Y]��Rٙ�5��;�@����g�V��`��M�MY�RVVy��F!�[�r�B���W�lZ����06�$'�yN��j|v�)5gx@�@�b��<�_�.8�ƛπ<9.49���VψCV=�x���"�;a�AS�Q���/�Bv�x�
��1�4S�<}xhG����b����j9�'����@���礖J5����i�� ]3Ţ�}QX^�\��k��;N@�5��P{����B 1ٶ<��Y.��
Yw�-��}ӆ"֚٫�I��7��'P5�r�2W+U��d_25gHt�~Q���eg�)�� b���h`��Y��?H��X���*��F+���y~(ܮl�DԷV�C,(	�0'%ۚntkP�mHC�5�Ics& �C��,�����Lw'��E�j�M�N�Ӓ 9��$G�C=�qz����ݱw��������]��Y�� ��.ܑ#b����%g�	�'�f}D9HKQaN�&��n�f$%D)�\�_��D�s��i+�yQ�ѭ�����;J��w��ߚu���?�����t��st��@p�l�͸+�ӱ�>w�Y^��h~������vy�%�6���z�?�j�:�	fW��t����@�I����i��h��
�jas���Ea�w�-u�R	{�y�!��K+�`c��x]"���,�!)4��*CA�{[;2�X�n�Pِ(�Z3΃H��-&���MNn�_�Bte>i�rE�:k'[��i�m<+�l ʠ�Z�i-��/o@�]!F����#!��:�,_�$��2q ���+�$��b��Q\�pa�௽�RnK�8�w��=$[-J�Ɍ~���Z�2�}���P�j����k�'�>�����n��KVK��?롶��~lO�<
~JT�a��${f^�?]D�������Чp�w�r`O�|�#ݡ@c�~I$ĉ��8RO;�}x�F�;k�ip�j�M���F2��������m�g?U�{�����Pʌ#X/�����ծ�.ASl�%��A(�.��p���"�r�4��R�w|�r,��������UyZ�J������Y�Ȱ��᭘S�T���־��z��M!{4Z���sˇ~VZo	0l&R��n3b�$frcu2�����#���w�W@�vx�ZE���9<*�.vI��p��:\�{�A�d����[��F�׮���*M7�ჾ#�MЖ��̐�b�=��LJ�����nt�O��I���{ϐ#�����Eo/w��5�l�2�5B"�?��L����B++�k@%�� C4�v�^*I�� ���-A&��32���'��oD�g��J��b��ף�޹q�?T���s���_�˓qj!dݎ������h�u���6��D���.��)�yBw졆�Ή��s]+�AU�ؘ�=��N\�/hR��0tG%l�m��p���?���VuH�i��حm1��D0Ե��> ��]u�Ka�{�@ф;+uΕ�L	pye�K�tG �t�\�4��^�ʜA5��ʈ�l#1�߆,Z!�y<�nb���ׂ���%Zy��X�!b�����B���4cJEQ�׍����v���%�~.hkC�Mꯖ��_�8�Ç:�I7�����=�P$���r�}��<+\����m�,`�"B�_�6ޢ��Qoih�J�40��t�����Ȏ���aX���a�e��ް���LhѼjR4b&�9�|�z�[#V,�<*f�q����!ͻ a���7��FPB~&V.�9����\�rYM�;��b�O�$$$F���|@C�)/a�@V3� ���!E���R�4%`�ڵ����-g�Ͼ%�����U�)cɩ��{����#�@�A�W���=�kGc��\x��Eز,��2y��(�����3��_�sn���fP# �_ZMz��;�u�_������/)�R�J3���($̘`>@�R�8�����D��Wm5���#c���`��yP۩��ƚ��'d�\3u��8��l Yѽ������S��	#�[E(�!<bg��A�u