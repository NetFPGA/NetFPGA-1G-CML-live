XlxV64EB    fa00    2b60���*~�-�F�;�d����fc��k=Y2�5�~�M�jz�p����;�I3�!�o�ӯ���~Yhs ��Z��_.���XA�L�c�����E'A��ۼ�[q���
a\�ȬR�bP��m0°���<�P/����v�ןz�;��hٞ)��z��������K4�G=ԙ�C�� �OR.����VٜX<�0���H*䡡.���{�/.��Afؖ�!�`�1O�H0a�RKP1���u�����]�.p����^(P�x����~d�p��i~��Å�|��`�C����[C#aa�<�k�lB��l�k5���z�Y ��Q[ۭH3�N��C��EG���\��SzaBq 0�+�� dƾ� �­9�W~+˘�Đ��?����
Q�7|A��X�d��?�	�1�/�0pG-,��^�� r F�ͭ(6U��D*�1��)Ȓ4$<f0����B)_IX�Y�ŋ�.�s�@�-�41riJj���qj�T`g�S����p�-/Oj����$�x8�snaEP�1e�RR����`�s��5F���5KWL�ălL:�X;D�P`(��	v�5;���^��n�����9c%��뻔� d,,�o�X䂠`ӷqq�!m y�t�P�V+��͕����`O���?���-b�8}���9&��������N��tR��� ���"�,ӆW�Fҙ�Ա ,uU>�I��e�<��/�*O���e?b�r%&�G�EmAX�I��J�Y^�Z�;ʆ�n`����o�ag���!Q6���������?�k
��7�S?c�r���1��Zm�
Ƀ�+���u��́q��軛=e���'�P�\P��ܙ.��.zQQ��x�^WN��~�O�A���-�ib�A)xX@U5�o��ʂ��j���sz�l7)O�߃
z�m�g�h���qJ�
�F�%%ҝ�+?�VW� ,�-xp����6y�AqU0��ǥ�+�?#�vxǭ�! �01�5����AR���6��b�7�b$�ȩ��W�wZRw��:JGL�]Y.�ޛCEK�!r���]�H7����ϾT��O��>κ�����>@7�ǔ�/�����6�b�m�ό�uX�oN�zT�3+����X����7z!�W�b���t� O�[�����^U�KY�D|B���g��a��Ͼ9f2���օ ��e�
Hl9H�?<o<�$�is��-Rnn�N�h� 9��gs��dZ���d�w�{s*�����p�5���O����n;v��!�w"�z�Tk�@�q���+�U�K�������<�B'���DQp�z9B��zJ�=B%v�Z[�j/�K����Q:.�t:�9���ΙA����;Xs�՞,�;�q�O=9x;��8ۑ��mMgU)�ˡ/qP\���±Q�9�kLx�.^�Ң7�U��~��Z�e6��}i>�U"W$}�c�ݢ0���\���-ۢcjlx�D"%��v\�:�� ZE5��fS��Yb�׹����s�_��.)��@SLX"�7"甡+J7���N_�9V=����QM`��\re�iZ�9�E��Bs�$��l�%Zw+h�I�����/����D%�5M�Ѩ��f�;���[=ٙhNo����W�Zi���Ġ�� E�Jh��ǬcI]��<|S�s�S)Eo+?�g�bRG~G��#�M���/��NȜ��� �&�F����c^�)u�˃�!�,3�U7Lgo,�!����vf,�뱇�\�h�0>P�4�G�_H	�@N��<�b|�IM%}��qz8`�A�|/���&�����c���`����.�ء�jM����~Z�$���R5� 5<R�)2�L���xn>���H>eIbD8�6�T{�P^!���r}^�?��MN���i�v���kѩ�ck�K<S��?�m	O��:{L�;�[|bQ폣`��ҕ�ݫe�B0��2>�`Z�����y��yZ�s�i����=���@����� WY�����Z-�r��#cMo���}���j,�7ץ����i[b����1�p�t��%��H��h��?�L���Sm�74Kc����S1qI8͸U�7�c�",e�c5Pw/6���W�2���kmr(H%�ڄ�K^�훾a��˳
�;c�Ñs�ݻ^�c'9C��؇�&G�����I�mF��	J��=�X�~w�6�p��Od�5�x�u����x?�:��TX�	���G�	���2`�����ٺm�� �)yC��3��N���A��X>S��(�M����k����<�
�*�r�LEI����Aљ^0���' ��
H{>!���V7CM�t��N|W���ߨ����5��_�Ed+Y�D`}��/T��oj7�&��e�O�T��V݅r�?z�]��-,jJ�A��P���<a�e��\�+l��ġ'{�n2��M-�X�k���I˞n��!�B�V۲�'/��	IO��T'�f��������˰o�꧑u���c�6Ș�C ��;�X�!h(h3�9��'�@˥�ǻS�Z�{4�t$���e�B۲1�H�k^�%�������i�dk�	�Ǐ/^cj�a��1	���M8]x�(�p1R@��������vf�,�Q�N����Y0t<�LԌ���p�Y�(��2�����~�W���w.2��q6U��4fS��di7Y�	��.��#��K0�D�֏B}�����t3�J
R�$��e�
����C�D)�B�SHq�Vm��ق�`��K� �*����TG�����͒g~�W��*k{��B��&b�D�AAo�AcsG�2G�{�(B,�t�I��y���?���l�W �a�aI/��?��.!m~#x��`	�1j��Y{��bTH~�!pn��@������2rE�u\-��88{B!�#KO�:<ZDڣaF��V����B�2u�JS H�M$�!�����E��S'J����;�ν��t	�Բ�G���H��s)�̤�c*,dy��Q��$�"�� ʺ�����v���j��?�
c�a�!~-{6���B�b�E�|���s���?�y��!w�X�z�ih�4��]y&��rG���7�*y��yJ�S�S2*���95h�#����"['AF8Hn�~�N�ZRQ:��,�n�~�D���a�0�.��m,�D��_��~���\��^���ޞ�e���#Y~����F��$#5����|�"�=�E&�&��(�C���� ��%e�a����$����H��zw� �at �QY<k^P���W{�X}��;u�o)�'�i����4MI��p�]���)B5�(>2B:���$�z�6�aEg6\M�Yi��`�	�� 8K����E�i�� �$�ӤF�G�F��,���^�ѿ+O��v�B@����D����񬉔|�v]p�ϔ�,��?�t\�	`ս�)�144��z�ha�4@�c�{r^����U��ǆr#����H���6S�.��M�'���Qkۓ��c���z��&�r�L"<7���'�N�E[�L�Iq?75�kw�����xP_`=�2n�i䧸�K�P����h�8'H|[�9�oa��\�X�s`%��Zu�$���m"���M/#�L��M͊��ܾ,_O��=�:}mq۲� ;����$ S��ype� �;f��d[����gb�b�(61���%P��)ڲp�z����#K��
���e�����U-�7��p�Ê�UJ� %�o�� ��f�����x�ё��Z�QќtR�gW���f�~!>��d�AC��_nKi?$�9��ğ�����t1u:������댄.�G�lAJ���֘�:�2 ���"����Q�%LW�g"�2�NT���[:H%P�� oQ�0i��|�D��������	��؅�dr;�����x����1���A�K}��">�<Ҋ�/�U�G�0��+�@���9�&���-���b�*���}�W�fGo��kB�N;Sc�L��&�X}O���R^�"g��`'�k��֯-��Bj��G]�bk���;�p�S�co�|g�����aT�U�l�:������ Ҝ�����j���Um3]��^�E���}� �MSt	H��=�\Em����G��W�d�~V�6�6���9�Ϯե/��C�K�GU:�CʬzT�Go�����*�Dv�`���c*.@���M��i����Y�Ʊ%V�X3=���fF ��!ح��Ş�|ƪ�f���]�*H��Q�.�
�|�1L���'6��+���ϗY8a��-��!�VQ�N� ���:��1��X�-ίn���=����}�/�p&�*��n(3�Ufu���b�'%�k�ƉK�|��Q����]4{��d��7h���ʌ�8n���@wV�M�Fw�D�nk�ȿlʂ�H�w*�#ĕ�W��W���fn�J��H &� �����J����NῄJ 4}D3y�y�&);
-�z.Y���D��/@.��l{�}�Ђ�#ǢBµ����9j���`f���|L��P�~��~��K�l���\�N
U��f��v��E����.7�4��ͯ}�&��z�k����1��qPrD<���a�U���#h�F��A��K���w�/)���*�5��o�G��2��J_����(�8�34p�G�{h�uVVMܙ������-N�w�ʯ�������}H��8t`�Smx�w�D�2M��<n�R��E^[�;R��ƿ��i�3l��G�j��(�p���]ȕN݃ =P\�yݒ*$dq~S[�p�Ǣw��ۙ%�>m�d㓄i!-	�Nr*KwͿb���A�|�z=�b=j~.�r��Q�L@L�T�}�����Ygq��T����!o�)"����2mJ��?����2�=��":��::TE�aZ�Z��+a>����Cp�7���[�z�	V"����<*D7>�t[��m��|�Q��t�jt�ɚV��G@����Cd�Vm@���S��{�4D�-y��#18Z�vޕ�=T1PR�.���JU�/,-s=�q����]\���8�x�1'I���>�i��=(�>g��Ⴔ6�&��g���8�h�Ygq2mu�s���[J�R�~b���q�vna�yq<�5�FC��A���H(Z�8����x�
���ߵy[\�}xW��4̖��kOv��4q/�Yj\B��}8��1��߂8��:K�V�`�^+f9n���X3ZH�A�@ڥ��,�L2�C����\�J��	h�1��Y�t7��)!}���7/������n����ӳ92T�ܢi�*�3�oBU��L?d���j�j!sn��癋;"��"�IQ�KU���(ty]�}]����x�)V�¿ �����ݲw�"�[������A3��J�oDӃC�B��R�t�d�C�"�Z??��'R�fn�㏂[|�Æ(���6b�ׁcߜg�:_�?�^��*�uY�[OLt���B>�)�k� ��A
�柪���EcS����~�uf|P�3D�|Z)���m�)'�	��;�,���Ǐ�@j;��]hC�E2��D�H6�X��h��M8��C�<C�[����o��^��	�;�3�4o�-{�o��/����s{�I*fca�rC���he�4P|Φ�5u�+śTOtW�~�x�?�騣p�,ro������m/៥O�m�R�\���;��Ő2f~I�-�'{��lq^���Y�78��>Q��|��~�����3-�18���f����Âk+1]������/�#Eyl�7 �����<k��Tux�/��^E6�	,ާ��yzR4R�����I�'��@f=��#;��i�O�K���G�=t��BbUs�+��K8P+ʙ�����u�nA:N����P��ŧ۬��X��Q&r&���<%�����2��W�����^���bv�\<�-�@{N�V����5�J!�[�Z>Fy2zA�fc�O}��l�'���]IS�H����Ѐ�]���n��8;C@���c �->u:�oGM�ŭ��>�A	�ig>@u�*��ᮤ��:���Y_�j�U�=�5�q�K@�䠧7�OS ���5���"��Ȗ%�b�org����+��K(	CK?ڃ�\E3���Դ�]|��Y̓�.%�W�=����.���)xD#r��/1g��Ǽ���C�����A�C7�M$��m01��gt�B|�[��C�c����;��Low���E9p�7�>z�$~���!w���c�1ѿ+�Ft,�C�.P��}���?~p�Q���.����#�	��T���%yݲ�R��p��]��f�1�4��:�
����Gx��lɼ5�_U���s�f��s��k��DSz��41��D7B���RUq�З(���CLB�#�B��AP�y���bcP��U��(��X���1�8�,Sj��!�%N_�t\�|��]�^EsN�/�8�wQd�-�=P��4^�F�󷑺*�6���(�����z"��R1Ǔk�*�d#2Lz�Z'D�サ6�Yi�ss�:�(�܂
<jV�{�e������[e���͜#q5�����B	�h�ë�gvR#�[m�i4��up��D��m�ׅ�BB[+C=w��LW� 0ٹT�jҧ-^�b�����l�B����;�kA�
��6*�� �!  #:�"�)ҚybB���D�k������#�-�H&���d�O�5@Ш�}������G����t;��-�Q��׵�m"p� ���&��Ov�l���t,��&�j��.J-���H��d�̋�J�祍�[�����"�b��$o�Fګ��1�9V�M�^j)�`{d5�M��17��*P*~�:���~��]? �`j a	����'z������x(Ti��q�-��F��� (z�pv��Q�	�TE,u(ŉ]�r�j,�~��E��C�0�`��V͝U@�E<v.S��׮/�#�v���ˑ��ƫ^�p��e�h�,�.�ĥ.���+x�T;aJ�՛M�"$TD�HG�]Uc��lv�r��d쎊��_=0�k�/�yr��p/^]/�d�Y��nԯ�4�=�,HrҒ��f����\U;������x]���IV��a`�gn��;~�f�Dg���lWG� '��"���[h�x�&"��9���{-��#���pY��g�a�<q��7:p�"�ꑆ3�K�;��� �5�y��s�r���HT�1����|B9���^?�e0��������7���l�Rj�8���h�vB�9���+`ᇬ��c��Oh�8O}ۀnI����sS�k����*&�:Sd��z����"Y@p�7�a�g�hd���g���0�����2�x
�Ǎ溝��k��<ަ.�$aJJ�}������w�0�8���4۳9Ќek%���h�Q��J�?�	�~�J�αc/$O��t0��d��r���?�;!��u�ii�_��8�Zc�]�����!~_l;�'�6���5���+�<7���l��w�{%h�b��0tl�˷�d������3j���^���as�`���K���4!�;�Y+xEt0_,Ri௧��\�[�f:I;��J�r��0} I��P�;Y@W���
���'C8���G�.�	\0Jj����4�">�ߏ�5o��}
��-Y�ü���q�V��;�W�eؠ�MZ3.�n�*2��.�ʤ3qԝ���]�B�$N���]�t��l[�6X��6b~���(v��P�{�/���&�U�����B\��E+�ʂ_�wa�
�Zn�2,��o���8��s��>�!y�S"��3C)����WiLt�@�?��.��L��i�a��
���<9XE���F�`�}Ɗܮ�I�2�p	]�B<,k0|zA�݀$dԾ7��p)��Sz��`���Ҵ��ϡ_�ǌ���#�G����O�HE�s_��ƫ'\��%��<��d̼�5̵���p���`
�[R����Ϯ�&��#7Jd����老���>~Trh�QtQf��a���
���S����u<� �:�ёa����a�%x�l9��[��xm�ʔ��ҏ�w�	�㘮�7����O=&Ǉ.)�;-,p���V/�=MH#��=���?�}�{#lק�j��5�������}��.��@��N�^]g��(?]�@�ijg��@��	R�c0���Mp[,���f���Ӎ����j 0bpl�L~�.����R�Ï��_[a��/T�Bi����E@��7isrz�ET;�f�$�/����1?���:}��B���EB��2e��;��+F�u��]
B7փS��;w.J|e	!����4�k��,o�ak�c_���LP��]IZ �Z�%&>&��F�pL��_FŁbYn[��������Ȓ��5E��`
��+D��#� �*�(�]�*0ؙ>y�K}-�Z�#s�'q �8�(:�BX���e����k�8~!�%�Y7<,�"�X��Ӎ�]Z<a
M�8T@�o<l���9R�,z2 ���]/�罺?���D��8'�"w��bD��S9b��]aw>���̲<dj��^Xms(H̎.���yL݇�OH;F2��!#�:�?���M�D����f�*��F�l�Ʊ�vt^�7X���yp��K���Qs���MŇ�}���WĘ�6�\�
Ժ ������T6E��P<�t�G{���	"�{��=��o�=ICB-N"�����H(������V�݅�4�sB~>Fi��Ƀ��~�O��I��Y����m���J�]@|m�OV#��q��$  ���T�"RG��(�{�:��~N���9gH��U_I/i8K�h_�n(x��b�4�1��V�P��Xq��5��_�>~���pe�_ ����ĺ���74�;�Z;-<�VC~��T��0��WV.�ꁏd~��6*))��>��ت�I�U^4C�qb�P{/�-��8�-�S��&������m�fF��Bc�(�B�T����o�O�#
��T���pǟr��l[�]�*�a7v�y��Ps40���30���;�-�5I��3Z��R�=O�6�@�(�y*Y�ĄW`ԇ���V��M��T�	�%trR ��@�9#>���>pEa��y�_��O�[0�sxKLk�O:��L�cEW��E�74�Şi��ߒ4ɋ$<4
Wgz�1ǯ���1�Y��,ى��C���5�1����ޗr�p����j۽��i2`zD;O�?�N���]�5k��7U͢k�1�
GQ�q���o�t��gm/�.��b̑ʝЮ&gl��[�%�h�}��Ŵ��-���FD=T��Η�$�\7��TJ,�<*d@~o�:�tWrOp�2O��J����e�J�:�E�3�o;����}��]"��g7�C�r���UI���Awvz�;�ܑ�����w��:������Pf�*hM�!
Dmg|Z����3��Z�wh3��n� �KM��W��V�6��9���YHk��'�J���;m
 λ�%��v��Gt��g��Pj+cQ��Ը���������w���>�o��J����KD°N�:c�����U첱�ѫ[*�³����Zg��җ�%�%z�*���h�I|�wm��O�e���u�
�2c#zo���4����[k%}���&i��m;���ɪF����2����r�@�8zfI%�e+������(����<o}�b�`��#����39�.�L����zԡ�j���ȓ�p��.Œ� t�4��;�p�~�_>��ANB�L˵���.8\اm2-F�`���%Ow�$�H$ق���0��i%�*o��.�`c�%�3�P�,t@�͌�7\��!X5.�C�?���l�9��Jd�J��"�K �/&"�69�x��Ryl�m��y�s�E��~7�*��D9 d<{%�]��C{ʼ���"KF���s���:=�'�Ԙ>5i�%���N=ǂo��{M����:7���Pw��U���`�6����א=|�@Jk��#�V� $��'#��D�,� �롢���LZ��򨩉is�Ү׶�r��>%�ə��F #q�S_A��l��M<�
�F��ܕ'��)h�0�Ўǝ�tz.~7�w����PbZ�#Zl��<Rξ)0D�3�Ƣ��X� ��n�]�����ш�Ε��v�~���2;Qr�(L��}InD-i��$>�/���pZn�8ڈ�0��)�0�,����$%�J�(h��F-5?���S�}@�ԯ��AI��!aՎN���� ?�>�q.�*BA:���?�w�IL��1:wK�:�U�����U�g�+�܋�"�ė9<�{�z�*��/����7ò%P�j"�P�>%�7ǽөVDN;qq���u���4"�.]���f����کzĽ0�An�rlKP�~����J��|�M�Gt0�YD������j��(���f�<,�Ð�Cheda�:#]��A���2W�N�e���� t����H�!�B��ٍ_6	�i�"
%d_*��u�E\�,I�9��G_�ꤲ���b�o��Rf��B���v��Xr���/��t8�o�n�/h
d<���`9����o.�~r�s+ާo��&S��ONʕJ~�y��ꡁ���!5��x�����o���C��r�D�8�J�Հ� �ٳ߼L�Jf�G��ژS@P#�4ru��O-<�n�0v�c������]��zD���`)ݔ�DW>9�Z�2A��S{Y� g�n�{��Q�D9�W�Y5o��S{�,#]�6��W����W��� �WM7\�fت����L5O��Ǔ܄{"*�W�S�eS��x;$j�Ft���<�6~v�L�>D���%zj[�3,]���2I�K#��� ������x@]Ya����^�4�a��o~����FC	��%1ǬU:�:��&t7��A�:��u�'�</[a�P����Q�F9�ʌ$0�rZ-K�ݙy'�ӭ���Drl5�΄�Ղ��q�XlxV64EB    9106    1830���x["H�o���?Xl&*r#�Lk2WC��y� "���w�'�[SԜ|�5��(6��c^�8�K�Fh�����2��ؑnN�j���t^ZV�1J��P¬��[��m-�e�	��n�������c�,�s2�!YA���a����}I;�+c�C�}�^�����Nᤗ�s<��X������'�`�g�^A�3�ʳ�*��x��/x�����s�KW����v�akneڇ�޹��M���*l�P�� �.ډ�9"e�F�q0d�4�%��@MDU�����8ŏ�I�BIQ=)߶ѢU�Ά��v�7���w�Pϥvo�(��3)���x�����0a>��|�#;f������H����QW���F��Ĝ��K|뽫�o��]hW�sR���P)6�0=�Q��*����?�V^<CP�Ed�-;���˓:��)���D����n��6�}S3��?����a��È.�_89믛�S}�	�2�%���@�3�?�z��AN�l��ܨ�U��|�N$|�8�����!0ñ�JG���b���aL"��- �=��V���Etd �u��e��0�R����br���YW�Q�SҠQ��F��q	&S[���E��-*�WBY\��'	_�[!gY.���V�'y7r<!Q���l��:xTs�L'V�7;%�q��P'���2sm�o�dc-ί���9�:�/��q�¯q�A��N%F{F"�hW	��^��L�՗P8c�+=u8�0A��uaE��Ǳ��[	�>�
��v���	ژo��$h�\�]�R �i���a� ���F�􇩮M�y�/�VY���S��[��6�>k�}�o��02�Q�˻��m:���,�.X�ئN^�"��,M����3�6%�E��Ģ7�J	�t�]_�O��i��]�Q߮�⇄��eg�dyG{�.��*����q+6�xG���WF�$z�+1Ͼ����@]̉;}ʌ�K���j-.U}��Bx�u,b^K�GNu����a���O�-��Uw����(���cS���-�[���q�S=�����$0�Omۼ�Ɣ�*'���sp�$�0����V�����/Ly��u[3 ��l<�b�~t:��Z�N�ҍw���s���8��'������Ϥ�0X3�r:֓W-���8^6���vu'����Zp}��r*'yz�:QC-������o3V[��t��as%')���/	�� O*�y㹲Oքx�D�#C���d	����Y?���2Z^+JmG�W��96B����JSɧÁ�n�L$���M�$�z����7�@�*v�R�0)�,�a�,�ۗk_��l�|�cN�sz��{��\�%*ϋM#E�;3�>�yE���+��N-sABi��{�{9�a���li�A~w�Uo���T-</׬�<�7�b=Y��{�h���I�����B]L4��!?*��S��Y9��e��$�D`l��@��:����G���Hh�!͞�8��u����"<�F���Գ�Mi��*�<w���=�����Y�����
N2����ښ,���:c�P籪���e�PZ;,y֠��߃dr��Z�������v�Ե�����]����4:�R���%�\�O�@#/��+������ �X��cڴ�c�7�kؗ��o�qBo{��v�Z�\.n�n�,l>G�����F�t�1
�O=�:�\Vj�D���"FW���Pw��dּ�����*�[5�-�?�s\���ш|���	>�&�����=ۄ�����EyčC?����+;�W8N(۪��E�7=�;��G�8��P���Ml�WT���n�׸w�� �_����xz�kt�R�{޲�&!�u[�º�`(�P�L\���+XF�
]��:O!��/r����1^z�������xw��:	y3���Pn��^���qݕ:�<w�~�N��\�*Bwe�Xl�k=P>`>�� + ��ԑ<�,�Lx�{N�O\����E+ $�G��{g`�Zse��]��M��>��6�r5��P�8j�C�� �o���ز��b�[~|e���JYl�x~M{P� )��1�͗��Uu\�"�cwk�U�ʺ���m/^(cN�'��*3 �c���X�ɒ!S7@+{�?�}�N�_l4-"�g�� =d����N�d�o���'��h�e�P�uJ6{멧+7�<�~�#��ǵ,�(3Q0Y����3�����S�F�O��������,�.�AЀ��Hm��F)��-W�����L�u�+���#^D���i���P�7��֑��^���@��D��|	�p�f>��ȏVN��`%�|�t�Ϲ�:�_B�W�M�Y��I^�%�����~�_DJ��D'��ǿ��؆x��+�B��E�U�?a6��8��z~���"~�ժ�zW�e�o����W�v;K2���ٙ�i?�����h����n	8�˸PL�.}��s7}oMp�������� ̉���5��Tv��>�@�_���l��^�͕�H\
�"k��zr�K?�����@gKrږ�fj۾w���A���C�(�m�y��&���]���$�R��'��!t��Ed뻟R�de
yr�;�����Z��ʉ��|�nj�N����[��@��E�na�Ow��Z�0}�/���yo(�A1P�C�$.�a�sK�sIE���@���Nک:&�9��<���V��5�����y��`(�B^`���tQ[�� �X-�:y;��aͺ>5֬ZZ���,(�im:�wlW4�L���)�7��b��@m1S��-˝2��5O�'��z�->�F�\C
�
��}KJF�AE1���d�È���J�I�a����cT���6���dG��*�b��*���΀���)"a��HzL8s��5��B�IvIC2?��~\uW�$t��5���d<�"Xj%kۓܾ����Q�=cvl3�W]��O��&V�rV��g~D�@R��V�t��T\DI�ųR�bq6	m4�A���6�!�T��+w�u%O�V:~��C3&���V�أoF-M-���FD8�u�Ύ)�,xD�	餝������+^��!�5-����$�����/�{� �5�ZAEY*(s˔��$G&��ؒ�q�Ky<����j�D'�� 	��>� �U��䅜��ݰK�7 ���꼲b6]gZ���E��TZ�RrT��t4���V4*��w���|�L�P�FWFv~�]�B� �܉�$3���w7n`c��R+�?��U�1)K����ua�2���s�
�1��6AG֝M��3bL{�����7v���hH5bnh�����d81AF213��]�O� ���}2�U�(rk�Ouƙm��@�C������������G ��\��Y����n�~��,��f�Z�Yo������
��ɝ!��$U��_IH@�6 е����`J��h�h��j������⻂h�iZX~i�jQ���Z�/v�u�ՇU�o�̦kb6�����(1Dך��l@X��H�dmݳN�Ϯ�t�_nb�UO8(��<m#U��&2Uv��	�)}�搁�+F
�O�Y�u�H�eý.��u~�����I�[�0�`���#��R�+�[�@5bv��a�+y�W��a֋����E|�j�P����SM%E_��i����6|��tЋ@�-�q�5��S�fx�b��!�~u�I�D9��f����"�%���&[����ks |^��"�e��%�L��s�HUv���Td}�S�)�y���(Ĵ�6�vt06�!�F�K6'~��a��\y����Dx*�o�a�b��e0i,�Ы��p��]%K�ʢ���K�4>n�lh�������EZ_{��/��\6h�>f7I�qՓ��q�/%L����h4����-����s�R[Z�X(K�7�1�T�#���S+C��KQ$l-OH��?����l����]<���Pz�L%�(�*��)�aGS����;��.w�G��S�ߏ+����{d#���k��ޗ���{��!Ƿ��@��Q;��ȌU��NxLP5�#]Y��=��u��"�Gu��s7�1IH���=��2{�x<��ri,1;jDa�S�c\��w����XS�Y?�����!j���QѡPrv�)��|C� �as��́8D�lv,\CHk
�e8 ��\'a6���Ҝ��Y�·�k��5��=�:D�yn��Qݻ	����y�F����&"����r2��n[=����@����ȸ�v^֋�Cs�w���bN���"�� ��4��T��Z>�� /��uk�Y���p�����¡0�����|Z��`׬�6p����3"�"|qB,Ĳ)���Mx���
��	�w�]��#�N"�X�iF����O,��r��%��fe0�/�?�;ӱ�����r�s�(���r42�lC�a�93)1�'+��SD�us��-L�|8$�3�H�ݫwD?��
��p�����Me�b�TuUAI��@c셄�ix��Ū�����N �z�I��珗��Jd�?��9F���TAgeg""�s؃�4��<2��_)[�N&�fM*̝����~�?03�P��W(����lb8��9�?��G$�9���3�L}u�77e�{܉��=�wG)P�_���kt%����VFY[ĴM{�1wL������9��O��^�b�,�ʜ����k&���ue�Ȩ b&d�d�e����a�Mrb/���[]�	�y�ٳ�}�������
�K�9�L�IR��.��8���\������I"��u�)�ʹ� C���'�Ӡ4_�[ٖ��@�$~�9��E���X��f��%�����2�Vy�q�~�"�j�rOW<jJ4���������#�T|:�4�y�;+�J�3©�F��� ������TT��ͅ�����L�V��i�D5A0G�(�Z�i]I��k��p�.���9#���
��a����-!^g|���8�@E���R��p����}�7�΀��?��a��\R�.e�ѐ��Ryn���h*�o�u>� b��6��o=;6��4������D�P����u�/k�׋�}��<�B��}�M�V	���h�̈f�Q1���@��7^�����5�펀�3̚3q�:�Ď��?��� ���*7������g�BX�Dp�vps�O֑����Jnq'�&謨���"W�:J��2��!C!#��v9�.x�-��9iDA��4�Wj�l�S��RX�d析xQ�'��X�F	�y�1C�w��H�`���|�kw�	3,"��6���D�����>~(�63��)*�E���A>ɱ�7�)�.��8@�cdiĝo�i�M��c��[X��O�B�:ɣ���O�^�?��	�V3!"�c�(7�Z�-��W��<��_�>Z�<���u`B���Jy�c)�ѐ��A9p ���[Sn���V��^o^��a���HW��o����O< zi�\'e�Ժ�n����/�ǫ�t��4�;N����<=W��|�fݵ/��F��j6�Jeh�J�r���V�~y�m.���V�����Bd�V�Ӥ�q���3}��GJ�;�B/l������>Z���Iߚ�b��{�`(Jy�.o��˯�Q�������F��X�ƕT��.��
�>�>3�8LXdV��٘qEh��l؀������@.�{Z�1�Wp�")m�$��(�����	=�?�	�b�l�U|t�t�{�I�s���}��rO֙��j���ǅ�Lo�<�	^��wȒ���}\l��[Er0im����H��d��^S_����^|P�;%Hw�k��Q�A�? z1��i�f�*x�_�o=1VkKC#����� �������_Ӊ�����!��\Jsw�������Y�����} �����/�S��|nZ��.��H�uջQB�T�m��j���sT	����e3�v���F~3<~6����%�;���+U���!k�`u� �X!T�[j��*8�+������a:���S6#�1o�J