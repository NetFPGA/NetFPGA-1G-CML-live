XlxV64EB    4a13    1100����b^
o�tx�	��a_q���b���k�wq��_ڛ4a#�Pc?%1f�ٱ�H���h���6Vkڸ0���c)�)�E�a��x���:Ꮲ����HiT��$��{��실:oE���8R�}iv���INÍzT�Z���)��XC��f�g�]��aX�N�i&h/�ؘqBZ�k]d���+\��<�!�t9<9D���O��'����� ��N��h�� [6�^��:���̓������P�������e�����h;ݍ&o)g��*ࢭ`�4z�ĸM�λ����4��ۙ��椨�*sXJ�Q�E�m�pP[��#8c2�xviG�ɱ5�&�OyJx�*�o�DKamx[��
p�>a��p,ȝ���	@^�2!�\�J�3�֢|���4�$=7�*e�_"�,��^�S&�r�Q��C���L���]�^Ф�Cg3�� �&�o<e/��x�Lf˴�j��l�UX�����i�ȇ�H�Y��ѳW?u�X��ƭVj$G.hh��n����iر�P�!q�^ٜp���'Bw0#53<��Z`YF��$]� %_�j_d�b�
?K%��f�MG
��
�/Ф����ͥ��	�]ټ�U�C4P���J���K�s�=ڕUf'gqp��۩磑���w��'���b��Ɍ`~]����f���6�#}Ӕx2G��f�/�	��mGl�m%�q.�`Ҿ+��R�p�|w	g΍K	ݡ��L�R�,_�L��S�i}� �����J��z e6���j(���_�q���^#���d�$��\�i=��q��E������������r��$w�@�3��kÞ�.Fd�Ɗq?����,�O6V��L¼�l��z^,�T�P�Օ�R�̸;����
z�N�0ي��lm�ߐ��^˪-eT��X�v��T� ��2���T�y�p�^���1��K�AR���S�en��m����v�#��ڽ���͆}��(�w�XR�OzO��M�|	�E�9��`Dt�����YW�!���Ω���$�lϻk�w̰`�a z����͔N��&���b�|Nc6J��G=6�3yk2"P������gO���R�ߋf���\f#%r��-���*�7��͊��F�%O_ͭ֬�P����6ZQ���[��K�m�HEb0�,���^�� ����L��S��T��5�ʮ�C~H�&(8"��Eo�x�}�㝍���fAU�Vc��\�C7�!L����i�l>f?"}�����$G#^�2�;b�����]�l��(�3���4&>�]���$���1��Jg�w�P5)�c7�H��h��x���\;ڲr$�:Qp�C==Єf�l�zy����f��nk��^$H���ew�%
"���:M�_2( f���%s$1<S�Ly������>��s��.���|��R?��?��{E:��$�kCf��q`$'Pv�w�G�>o
{���2)�6��"ǩ�^����J}�D��<bsJ-���|��5x�+����v�z�*��8��&%z��p�͟/�z��-����ե�1��Fg����'�y��8-�����T�pD%Z��R���b�&{|��T�)>�:,��ծ�c��o\����H:��o�/-wN��2����L��됪��Q�_�'�u_J-	L��$n8�7��TM������d��}^���������[-t"J�z�ssi²ZW,>B4�o�}]��clM����ۋ^1�ǣZ~r�?)�Ɩ)��.2z��5I�*{]o�܀�d�[WY#����?�z��Ɣc'd���HǢw��,���JI�`�eC��0Sɉ#���P�Y�8_pU� T�;	���n˥>��@b(]��n�"�@!���M`�kWJ�WD�>�Z�[q(�
j� 
f�2tF7���6�w'�$��t0��qG��):��s��ǧ�q߫��*�h�gp�+s
�1��Iaf8?����n����[�%��ʀ\V8��~��s3s#���@���<���C�ʪj-O�	#��Ý�`�����֢�c6]���x�Ն��TY�|y�@�f�O?0�����K�|�4#�aLhMՏ��k�p�;�v��8�[a|U
hl��6�#�)��$O\�y*��^����da��[>�6��r�kiY%=8��P��~4h>E���N3�����O^�F'�%��v,>3Ϻ��C�oɡr���+Y���{���b����:�NH��I��m ��n��W�Z�*��8n�}&���|J�+HM�E�6�Q{
Hx	������:�a�7$�j���I�w9Qa�\�l�&u4�9 ��G���%�fώ�	V5E4�GH�k���e#
񅙍���1���N�'E"m16zx�>�r��=��(ƣ����r]H�E���g��j�q�� ��cZ	\��K=X:���*��-;���I��$|���I�_�ᎋUt��?6c)�͟[�J�S�il"��{ĥP�G�@��72icd;g��� ���F�U�nu2��)U5#|vbO#?�AU�/�9��k�؀�K�R�,�@�b�>�c(�%^�{R)b[J虷|(8k��MU��S6wl-5� &������Y�.�s�,��w��P���:�zd��%*�*M����$��j����ɯ�8��V���`���Sj@�M�V<�d�P����k�ly��?(�X 9�n!=+�D8�ͰR)���IHD������:�ȧ�X�p�A���������D��2��i���mu��"q���y)�Y����5�R*��ph/����U\�6o��M`�x���[��c�`������k���BXD9	�����:	_�˷�g��O�����Tm|:�ne��a�������@������ޠ�3��U�'�0��eay#��iU4������粂&�\'[�z��Y,��{Y�j���2Zoz�J��:��i5���(&Z�#M|'a+Y1`�W���-a}N�Ȟ��� H�űOt���!��h�u��(��ֆ�9LNp�F�Fc�:�����j�t�;���a$�u�����Y䨝�NoѨ��s�a��F��O�&X����0��'^��:`����,�Y�Kp%�M|��P�ʁ]�mp#��(�����߸� ��������N�-�#x�A��8�0$�|#�� �Ϝ�+��.��Fz��v��*b��H�D�y��.n$�K\�^��&���ӕN'&"�PF�_:x�!FC��ش'���0sF�S���~㛭��+���_.	�c��쓪.�kxx�I��"`��j4f�$���w+�u�\���� -���~y�-�5c�|��������W	�%�+H�M��t�_�$���wk�+�`��U��6t��c`9	8��,�6�*p�;�^���ibx1�"�@fh\����أ�����m
�A�Z���ζ�'R�cĮ+"��x�WЛF��\�~��s���֩��K9'���Y.���3�Z"Y�[{4?{t�>zjG�_����˂]�	a2�^H���9�Sh�"5����-J�Ť6��d7�^#m҇*F���l��htI	����V��l�� ���_�E�/��愃�جԠב@����
3����H�&�E�(f�ߛ��h��`�.˙�����ͭ ��!@E�T`�fx9eyL�2�o��m����ؚ�{�tN�����3�^"6��#h=2�1`Jh1�4u��\[Hզ�f}�2f̣�I����8U.���L�W{�mF~{��e ����/
�_�f>��(R�u���𞣄���IyՁdl�y� e4���]d<{��͗�1���*ƂE�#Gn;��j��d�:^%�B�ڠD˘$�.���j�}��Z�,H.���|Vb�s��Ӊ@^�i�93=�z,\�x��2����8`�g�-�cd'��ah[���m���h���=�Z��>�d�K��� ".�e����
��~���/��hR���u������1,�DҪVy����	�n����ud�_��0��T+	5�3�
���x
��:N��){1���2��W����g�+
���N8���`4�?�&�+���#%�s�L�3<V���tj��[Q}�Q�%����/�8B�� *ڱke'l�ZnU	 I��)^L;*��^�X%��Ow�!'I��Τ�S��
8��_���w;�����D��s���%��_Srڌ8׻i�%��[�IE '��a:��0%>uٟV�[J�����6,��u4���