XlxV64EB    54cc    1000[�
����
�0���8�Z�=y�\���G<w���SC�=71(�6�@����Z�b�g����`�fc�>ȣ��z8���?9� �~F�P�������<�Q�fra��ف9��&�e����p������Xt�y���4��U0_��^�6�Sp	2b�{���dqX^=w�/��8��p�$,���V����E\@�B�V7.����{i��D���i��YS`g�$�$.��>�ZyJ[�.���.�Q�C\;+��а���<P�%T)772dl���x�gӡ�����@���V�MG]����p�J���Ʌ�:u5�V�<.v�j��:L��5��u�|�@�#"|B��6��� ~��@����[�1D�^)E9�o�Ēǎ5[D���\H>M��>�iv7/}��F�j�ي���U\�L�(0:W��fF�RЧ��⃱d��A��UQ)���E¬��~��q�T\9�y܌/�~Q��������exL� 2�C3��>��1?Ut7�@#�7�f��ǻ"�][�x�8�	�,��6䎔����&��`�����:�%u�����G"����@ `2���yf�B4A��e/��u�6��j4ш#EC���գ��$�KVz�+�&x�m"$��p��y��]g�O�����C��h�Q����VH���Mb�q�A[g=�ܴ��5O#P�M�6|�=�T!�����
�4�Y�����𑮌y�aH��M�w�W�)�6J��J"fێ��ܿ�z1�C�P�$q��l� ōb�P��A�����B� Pw�^�Cj�`��E�"�[���d˳�ށ?���C��߇��U�m�f�+��εs�y�u��B����,,pP�֛|Ay�i�-@���єYU�}=�P���e�GN�F� �!��x����AdvL�'�E���&B���!T�=v�� ��|N(Q,B͌uKh2˭ ��ZQ���/n���H��-~2rR��m���I�1��y�8��,����k�*������7Ã�@u�2��V�,*"^���
�ږ�V[�����U�ZzS�[�%�ڄ�� �4���h>`#�9a큱6Y�+eR������h(P��ZN����/�����Tv�█�~�4�Q�\-������{S�Ԯ ��33�D�4�ܠ`��Zpڑqв��d�hy��pG<��_Z�>ғ���έ[˂�>����� �r����g���$��h۵\���l2��_D���A8�~d��2����R�[��7��E��z�_�XIj"a�[ a��)1�Gma�Lߘ�G�3��|��2�c��� �'u����Ϙ�ڞq�?|Mi�h�&�����=��LK���j�ȟ���-I
�6�_���xJ�G��^1ڞ�����w�:Mw�R6��%��.���n����J��<��Ίy d�K�~2L������)&�:��qHY�ح�XR�ҵ�?0����k8���H�8�n�H�� k��8�~k� ��rkKHl������L��Ǳ,�W���cEG�ƁG�v�ʒ;��UG�ą�z ��V��5�g,ש���}���6d���S����j/�5"�C�l�|�����/k�l�5J�9����4ܡ:�/��Sb�r���׆�rI%�YA<�3}���;	�HS[Q�G%�����g�"Y>�?6���*����@��H2� �^o��R���N؆&�0H1X�Nt����5�P���	��Ȭ?8�Yo&:pVo������i��6�5���m�9�hƸ
�K6"��]I�GJ��>�Ӵ>_p..�s��� y ��2.TN�Ӡ�U�c�d���6��(")�%�LO�2�*k�f8e�㒆)�hE�� bK�f<� ��e�z�Z�,�|R����In��LxE��KcJn`�O%ǻ!1���{$!�C�^�N��2���y#9L��!�0l<���$Ŋ����iT�����?�ૣ��:3����% ˴;�(���}i����߀*���`6s�����pvR�O�/뼮Q�ᕰ%g����ǌ�j��8B����!�d撝���M���y�49'N�8r��?t�l/>�c���F���ȉk�C]��6�)%/딕$��j�ES�]ЇS�{�Ծ=������X఍�{��l/l�M�?;r_�t�Y-E=LF�8}]�Me�m���}n�����5����]au���SXaS�T�;CF�������Z|z�����br�qSsgϏ�e�4�>��	v�%�����gd�d�(Y�埗�c���3�j�� uB"
�&)�P�p]�ȗ��cjY]�lx/%�H�*�U%Av��3����M#De�=*��*����0�v��k�?��\�2�9�T�b�=��\]��_��#�����2]�~��n���~:���nF[��c�5]K�	a�o��6��P3_9��p�~B��<�A(ʡ*2MBV{,���~��W�_ 7=4�q e��,[�i���Ƶ���7�[�4�Ѐ�w�I|56js/mC�c�اKq
�J��pv�s���[��ZH�gO�[�BjW�:F��]�6��ƊhE�P,����7�R&���V�N�הjQrg.��&�f�I]GE�lv�sou�/�;�jv�Ӣ��]�t'��CZ��9�B0��9�hm�T?��������Am�Q���iY��a��;>��Hf|(c��E<�Ht&�{o�\�֌R(���V��ąa�� =�բ�N�u��o-���ㅃt����?h���is��ə�Γ��+�I�ӎ�zB��n�3?#G��K���5�O�����6/�R��<x�w����h75��l�h% J����X�7v\������'���{f@���S���r�Ѻ-&�<��qs�2TG�c�8QХ֡�bU�K�}_׊GgՈ�Օ�cz;g�h[�ӊAV��޺�,\|�ʘ�W%-#�Oo*%�L)�5�����!��#�9����kl�n�]+��>�<���L�!}�QV:G f����-���w�CJ1)����ܟN�Vv+�v��Xjz�^���8=Y6>�Mjj�k����ƿ�$JO��ܫ�QA�\.y#�YG��'�.T�Ȃ�"���3M
dV�+9]��'��Hݖ��N7�n�<}~G�����kWS�h������3�V2ۚ
���4��~��a�o/x��c���o.��C��F�E���,E_c�����7Z�i~�������v���U&O��	��+BD��V��`��4�K ��ǥ�l��l������3_y�/�r݌	 �R�"�@�B-EM)<���> �XG� u���v�(!5d�Z��ѶXJ��7)}�ٹ�qIoa߄��X�8�+��X1� V�_68;x?�>��w�ɣ�Ь���u�loO�������ֵ��\o�-˹��c��C��8֩�ATvW+TB�^�����ei�.H)xG�2�.��2�`^`�Dy�^�/b8�I�9.*)ݴ�����\�����LS˹foJ����T�꫆˚1N{�3�эȴ�e�j$�7����{_���QǇ7��X)	A���MX#���4��G����ǋA?�c�I�������z-z����X\�tu]���lF��A�o��Oĸ��9Rh��6WJ�pe��(�������/���:����6x�7�Y38��ûR�%�00����!��݆�vS�n��z\��S�(��3���E�V�@�%[:�����[+���[�ĺ0� ����L�����xop�~ȶO�I:5B��=�n.Ɇ�Z�6��ģ0�r�m�$�;�@ּ?TU�7&�� ���D�t�F�����H��`N��������b�o]�=A� x�\���Q@�ƿ�v��( e3�Q��]��6�z�[J��<��~���d
;6(����WVM�lw�����=�¯E��~X��CVL#3!1��D�~-e�V�u,>>�}H�� �Es�
{K3����ٙ�bX�9�-=���g�2Ұ`���H�~*��OG9�QB}�?��A"27�+8i��Z���o���=