XlxV64EB    4110     dd0v�6�
�6��B~7���[`�.z������ �ylp>d��v��Fݳ�<�j�_�ХL��n�8fu�ך@��ʐ� �Q)S(|R\H�+��O�d���@����d}���>u�wܬ�
�`��DӁm���}��;��,�*cɵj
�_�2�3mh%٘��.�m[G:Eʹq�"y�W�5�I�?".�q"�x�#���� �ҟc�U`�ʔ�����!L`������_
�	��pDw�+��)�AI�(��-��[�s"�r � �)"4�xSm��ΗH�ژ�ZYI��^+�8Π�����hG(<Gq�r�]G4�4 q�C�hhA�"̗�� &��ք(�Z�L&�߳5k攽�"�	-��_vf������Pbwa�-�J��sf��i�Q+�����D�)�kVɯ�����pC�W"b,����~��&4-��W&f�u26z@���:Dر4/�Q�ԟdl�`dv�jˑ�#�����	�&yI�&�Nv�C��*�*��)kgRSj����=��pj\�Z|Nӫ��A�3��R�D�<�0iL��6Ё�5��`���0�j;hUN��ԫi���r�Ek���-&�5��ùo�W
��b~�ʨWw�n�JQ��͛o��	���oe�{^t��;��"�����`��B�s�s�B�^6�C�@ơ->�n���kc0� �AV���x���_��@�}0U:��$�ciD��l�EO����9�Kd �!�p0��Z�-`�F�u��e�,��`ܬ�e��퓚
j#����՘��BL�����{���j�P*���a=�s��Q�1��������9R�b�N����-���%*���FgS��ɜc	�E�/uڬ�u��8��Y���0�OnA����4'P���'T��B.�f���U_��G\��,,0߆$&�Ho)Է�/�r�����w(�v4����BRO��m�XD����^U���o��#����N~+�ʝӉO�k��k�g���e�'�vb�/�N���B���JN�m��[?O-�v���y6y�.u�)�[�	�E.�c!�ϊ�D�R���U�%dH���j!�J��!�_�����vN��Ι&-O*$�N����#X9B)�;��Y�o*N�C�>͑��%_䢸��j,�0}��a�/c3g��9��@�pT��j�@���^��x�G~dq���p�T��ʖ5y�˼<QϮA|����l*�����_%���b"���%M67��zx�􊁡1�>��(M�؝�L���S\.���>�]�|�D��Y.��70Ub�[�/B~��_l�;e۪��=���`����:_��
��ɺ%��UD�.�z&����Y�0��%nq�H|�D���u�E^�_^(C�Gm�]�a�]��)#n`}ы����l��\�{l1�{	��/��zb�El��Im�����~�x)�Φ��{���,m�U0*�d�B��w&�x9-к���R�W���1�S>�&��mGX��!�D'�g�&��<m��R�|�n�!Z$����䱮C�qD�4,S���a��u��w�2��E#�o�ޮ�t`H��5U�X��>����| �A5�ՠ�����Z�P��a�S�2��K�ߞ�zC�$(�]Fw�Ũ[7�u�h�~��+t�)�m���5�	gҼ�,�f�&a���&ç�ʧ�]E���̫ԟV��ι�:���t�6l�5�	#Y8���;3�W�ǄJ�˘&.�A���>�W���R3�/�*eYoL1����{D��ۑiG(U"�jW]�%Dj���E��&PA-S�:N=0͇&�Lu#�8q���R������1&[�E�-s��t��r��e�ڎ�������K�ҀިSc�L�\�J3 ���0Y0B�b��bP��
GU�o=����N�ula���,	W��'G��W�r�7��
��.u��m��?5��}�'��1���r�*��ʙ��W	�cS�։9F��>�i[�Ql�&<����a{7
<��-cV�r�f��z��0 ��E������п���/:�Y�g�K������H�|�&�O�NA��Q�z�����*qH�`U�Y<]6B��B�Wb�aӂ��	�d�K��\7�g�F�N;3ߪݭ��e�f=�p���f�!�g���ֽ�<'Ql�>ެȔ�#�Lu{ʶ�N��vU�8�o�QW0��*�0e�VM_�cm��]Ĕ���%�C�+6LG�O�R
	��C��{�K��6�G�E� g��W�#��P���v�Q
2�K>�T*+	I�4������ȵ	���ּ�V���SX�	� ��
��+6�����N�Cg9S�h�	���V�p��l�����b/v)Xe�P?�����P�U	ŧ+�K�<��0U>oW�-� �Ҫ'�~͞i����3��1��P FoRdR���*֒�CY?�N����,2u��y�{���#~�n�H}|^3:T���gw�%�6����7~E`�����)��e�<��
�pD%�*�yc=b����ب�t��}��ۇ����˵�5�I�:��İ�6ꤡf��P�c�2���)�^�Hs�bB�5l���q4�{�^Cr?^@ ����</��	|��	�1(��Y/���-;#S�d�3��d�w�d#�52� ֭�E���y%��G�4%�+���I���آ;ͧ�����W����Rh.��E۹�Ō�0#>y �Pv��9z�fx�9����n�&mb����Y$-�O�����j*B�}��%�V���uW�+=ߴiL�:�E��{y?���aA{x[1a�o)�W)�q	���ia��[��)7����̆�`�����k���Ǹ\\���8���Qt��K_aǬ�#&�_PHoB6�aT�-��V��wEt�L�ȭ+��8*�7�'�,�8�^Ċ����������lN�\{2�[n� s���vq+��;���dK�3.�ah�3�i�	�0��+"e�ML"�JHO_�֏'�^+%��;}l-������	Q<���]���ܫ��s	ɘ B��W[;��%5u4�z�g�h��ŊE^Z�4Z۠��_Q��F���l�ƒ5f�~��	�:
Q��)��"���r�1�}�_�S(q�`��}��Iɥ<�u��5���Ġ�؛�_4�Z�d��TF!���k��2������[W� N��ȷV6N�s��k1%G�
bg���q?TY���[,���Q��W�%�Mn���&���#[�5�tf,M�h
RJbO�HjFWN�x�?˭�m�z��2OG�lkOɶ�[��q�X��r�3՛��*B����J��ʘN��[�Y�9^��t��$��{�����O����ŚKnZ����P�r�߶:G�y�;�u���N�%܃�d_��P�`����.Z�D��:zxA�ھ�!Nۓ����b�CR���|��]�zz����K3J��U]KN@�� ���<��յ�4j1�