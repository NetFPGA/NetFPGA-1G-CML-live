XlxV64EB    59d3    1410��j�W/5�a܄U㣉"ا��='s&�E�
`�j�����t�,�+����U�mld�Rm'�l�SѠ^Hl0WN ���-!;�A�z�Nt�w�g�S{�g��7���K�ᶇ��X'�m9�����i΢Z(>�8l9p/tҺ<���6��D�������|.�������^p+���p�I{b�WC�-q����M��l#� ��՗���h���VI��0ۇ�oX<�6��3�{m$�G��J;�1v�r/��Q��� ����҂!�!)6B@��-�3�PS}�t�����I̝TG���o(�|�7F�����Os����i~�h�|�O����*L�S�9��R��h����IW
�5�������?~l8i�<��Ro����iv(�2H�y=�V��Z�������@ۛ�Eg�3��ř�ލ�1������*�����9�������N��_��Q�I��OBD�\FF�~�惍�kaD-UyĘvʡ�hTB�
���y�2A*[_�S�w�ι��4�"�_�i���s_��+�FP���54����m�P�������v�̨}��E:���ť��<�8!`�z�{�N����2�!L̡�S� w�e���#ĺ}z����u��k��|#*9��DE��0��QI\��E�y�e%ի�u�8 �e��#���l�����K���x��Jl��e�Ri!���,��1���Y����B>�@1���Q��ѯ�8�0%|����AI���HE�y��U?��#��oW�jI�Ip�s&}- ����,�5�����J'p-�*ǃu�έFH5�)&��t�*⌲��1F.�7�$xME��ͥׅ��jl ��^�+]㯞�e�K�X|S��NUE����c4X�9�� �z�����PZ�w����7����g�b�T��/���uO#�m5������ c��\7#�$���������[�cQc��𽻴T���!8�T�"V3�u������#�kA�>~� U_�.#Z�Z�P���5��2� ����g�`�Jq5G��[���}��@&gՉmp���bڕ*	R������Í2*0�N�`�����M�{g������������\%s����	�F
*c$���3��N[r��w���tΙ��m��4g�����Qι�#A`���F������R�G�LсZ;���l�g�;�t+Zf��3��X�����&�̱�"5�+����4�5�,��xs.��և�C￴F2�JL��?'���D��}��1 wx(ϋ�x�@����h��0�A^0�������;s�ѕ]��5R���΂��vz���n��m�ҕ�4th��0%���kr��쉻�MJ�@M�QU������9���Xiq�q+�$?&�����n�s�0��F�{b�w���ʆ@�陼ɷf�2�fx��b�Rֆ����c���	ߙ[n�I���E��i�Ӊ#���]�ſb�~z�m*��I-k� .`�� �����G�E�P��X�@)f��U��B�7V;7�nb������E�;}�Jo�o�~R{��^t��0��7�t�F���r@�w��b%؁��$c�$(V�;s$&�8�$��B��p�v��h{@/���L�U�~w:Ӂ���4	GD�N�f�ݽ�����>��K��Y�O�ra#|��B��Ϙ�4q��l�N�����u6���[_��b<Pi������	�G%64��\C]0��rC���z�G��w��Ҫ�2�xsUxcA57�Z��&��>#���Ȼw�`��j��j��6��(�r�]���!�]��3Т�i#	>�_�i���Q����Ѱ��q���yV��6W�_��?�dh���Y<��+9�M[e��A�eu���E�Pfr��4�ɘ
���F	��,y��QD��xC�(?�I�6����N
G+�7�[�QC�?D��^� ���44FF+5ےn�I��<������M���:^FY�Xb��i��(bX��&e�(\�e#IS������QK�;��u����.
��j�ōX�4��!�0�����U�����JYBw�tյ<�y�&���t�/�>��,,��{;��rW�:̠99�4��Λ(|�,���쏵zwYb����F>��L�e��וk��wn�W�K�]�1�Xr����ȞO�?\�4��~�r@��'���Yd�@h�9��W-��K�`���'jL���U��a)�������8�񱥖�Ѻs��d��l�4.D���J����l��5�F����N��{���~Y��(�H����VLx����E&5`�3�#��m[l���^%^?�p��{�46������F^1� ϑ��3$򠞸�55���G�$5r�Y��P0�w���)�,��F���m	`+\���w*SX�j�
Cr�T�X��x���r��MR�ŠC.C5m>��~��:äCm��h����WC�1�E�f���2��c�O\��? ��U]���2qk� ��cA��/o^�<�ـV��_&�}�ZK�1�?�$DjI���ƃ5TD��h�ϟq�m���/���9�4�E�z{�ڛ0U�FN^)d�C�}��*�u�y��ȋ7Xv�X>�!��S^F4Q�Pn,l��H���h�T���ƌ��U9�j�� �����Ј��75rW����c�!�eG!|�������$S���{����S��<E��!�3_Ȱ���hg$y�9B�Z4^T?�vH�o9L������]�S�T�Q&��\>�j
/}3�eyC��J�p�)�x*�_Ɠ�� 7q9`��F�Tt��U��I��&���z�i��.ӊ����U\QK�D�����e�x�<l*ö�-& q��늎����7�� �V^�UQ9�[��v��Q�
���J�PY���A�~���S/��Ѵ4m�La��6����f�i�u��}��Y��\���+㼲��%6��F� �b����(��Z���n��L�k�݁��!�i:�/���"+�l��J>�x�PJt�\��ˢz ��e�9Hөo�����},|"����ɐ/[��Z�aA�{�	�s��Pz�鴨,5�l�+�����rp �(*A��!�>��ӞC��>Oo(����B"��,����f�wf�3��p��Cڪ�SK�0�-Ď�+W����'\���7} ���S�Tu�5�R��f{;��(�;� �r��8���>ʖ4��,��nvX^��fRv��<��kc3m�`+�g��j"��2�🮅��fq�ͪC�r�����b�mw��Q�|���!�s>�� �� ��Ԅa_���'D�t+���7I̊?rF����bA�Aܧ|:nr���is���9	|�s�ڨ�i�S}HD�����,WOfQ5�c
H��4 I1�W�F�f,������l �ڢ2�aiB02�zO�C)sA��=< <�Y%�0�����j%�'vM�Un4-y!�]]���[dL����M���񿼝|k�����Ɋ�ԫ�i���*��H�o(�Q�Q�^��6�s�M��M2�GAo��^�2ﮦ�ڬQ)�=c\O��l	^�=�B��31dvq���+FV���+�E��먾 ��F3h.Bmx�x]��3�}7tB�:��!w���<�cP�I��\�M�������e,��%-��AT��cػI�Ϳ���F5<�>_?'a��C1�ʊ�n�y�C��+��?��B9������;��N"�f%�8�+�ܳ�[��߱\��{���ܡ2�����OP�o^.Z��,��N��m��)�1 QL<2�sjpd�6�<�r�Aڠ��B��l/��7S;�g�+}1<m97(Ȼ�Vר9�m�
���dJT�*}�;��.H��9K��J�qWp��s�$���	 ���O�<|)T��T�A`]ʻ��?Pg������_$�F�J��rP��O���!���q.�*n��%�Os�t����&��")9����>��8
�n73J^����Z�o|5o���'n��P�ɮA[�.5T���G��>�u�0�-����7R�����^���k\��aw��S���-�^�V�l6���L���Q�Ϥ����w�!�՗�6-�)%f��`޶�ڗ���������m���׾�Ӂʜ�X�Q����@�B>(S���kXf�1-G�'�˃4çD턈!�Za�q'��~�������2����Ν�k�8�ќ��!)�d�/�-��/��b���H��w�˲��[L�x�1� ;.�{��$�Ѯ^p���w���
��Jh�X�J���kCO�����j{��"� ��*B�`��E��7'7K�$�mGu��?�7�G��	��	��|��X?~U�������Z�F|�c�*���o���`�{��\KJF���7�wG�7����s#�chQb�̖l��1,��8��L�@�z���n�k����[�HM���ib���9Ӽj��̀�g>��'K��|�L��Մ^�e�l��m�g#[qWr�M�cX~��Kp��G�>3��h��>�:��p�E��2�tK��D�(�[��:�8L_�,"�{�j2$�G��N�Y����"��s�>��W�?�q$��R[���+T��`�[D�DK��?'\�� h5��;�__�Ya�c��r3H�����n��ħd����[h[	b���%
�wsD��9�4����RVrDay�3��1-v�ȅjV�0vz���,c:�bư\�#��8%�:���� �B�(��_6��!�R9�`�b��5�}�̈��+.œn��(��Ҽ7�}h�����V�Ͱ$Q� ���7�{B65;��������U�_�)U��8����D�Sv�ߊ�ax��Ts��%2>ejӸB����NIp��N��w�毾qpJ1+@�8I�8=�U��⺤���st n�F5k�_g"C��W�7eb���s�q�@	q+�+Z��md���u�I�}�����#)G�#<x��G�Y��h��&W|&�C�Y���Q�A?iL�U��,��8�Z0