/*******************************************************************************
 *
 *  NetFPGA-10G http://www.netfpga.org
 *
 *  File:
 *        cpu_sync.v
 *
 *  Library:
 *        std/pcores/nf10_regs_common_v1_00_a
 *
 *  Module:
 *        cpu_sync
 *
 *  Author:
 *        Noa Zilberman
 *
 *  Description:
 *        This file is automatically generated with the registers towards the CPU/Software
 *        and is responsible for clocks synchronization
 *
 *  Copyright notice:
 *        Copyright (C) 2013 University of Cambridge
 *
 *  Licence:
 *        This file is part of the NetFPGA 10G development base package.
 *
 *        This file is free code: you can redistribute it and/or modify it under
 *        the terms of the GNU Lesser General Public License version 2.1 as
 *        published by the Free Software Foundation.
 *
 *        This package is distributed in the hope that it will be useful, but
 *        WITHOUT ANY WARRANTY; without even the implied warranty of
 *        MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
 *        Lesser General Public License for more details.
 *
 *        You should have received a copy of the GNU Lesser General Public
 *        License along with the NetFPGA source package.  If not, see
 *        http://www.gnu.org/licenses/.
 *
 */
 


module cpu_sync 
#(
    parameter C_S_AXI_DATA_WIDTH    = 32,          
    parameter C_S_AXI_ADDR_WIDTH    = 32         
  )
(
    //ip clock domain
    input      clk,
    input      resetn,

    output  [C_S_AXI_ADDR_WIDTH-1 : 0]             bus2ip_addr_sync,
    output  [0:0]                                  bus2ip_cs_sync,
    output                                         bus2ip_rnw_sync,
    output  [C_S_AXI_DATA_WIDTH-1 : 0]             bus2ip_data_sync,
    output  [C_S_AXI_DATA_WIDTH/8-1 : 0]           bus2ip_be_sync,
	 output                                         bus2ip_sync_valid,
    input   [C_S_AXI_DATA_WIDTH-1 : 0]             ip2bus_data_sync,
    input                                          ip2bus_rdack_sync,
    input                                          ip2bus_wrack_sync,
    input                                          ip2bus_error_sync,
    
    //axi clock domain
    input                                             Bus2IP_Clk,
    input                                             Bus2IP_Resetn,

    input      [C_S_AXI_ADDR_WIDTH-1 : 0]             Bus2IP_Addr,
    input      [0:0]                                  Bus2IP_CS,
    input                                             Bus2IP_RNW,
    input      [C_S_AXI_DATA_WIDTH-1 : 0]             Bus2IP_Data,
    input      [C_S_AXI_DATA_WIDTH/8-1 : 0]           Bus2IP_BE,
    output reg [C_S_AXI_DATA_WIDTH-1 : 0]             IP2Bus_Data,
    output reg                                        IP2Bus_RdAck,
    output reg                                        IP2Bus_WrAck,
    output reg                                        IP2Bus_Error

);


  //Wires and signals

    wire [C_S_AXI_DATA_WIDTH-1 : 0]           sync_IP2Bus_Data;
    wire                                      sync_IP2Bus_RdAck;
    wire                                      sync_IP2Bus_WrAck;
    wire                                      sync_IP2Bus_Error;

    wire                                      bus2ip_fifo_empty;
    wire                                      bus2ip_fifo_almost_full;
    wire                                      ip2bus_fifo_empty;
    wire                                      ip2bus_fifo_almost_full;

    wire ack_event;
    reg ack_event_d;
    reg ack_event_d2;

     wire read_en_bus2ip;
     wire read_en_ip2bus;
     //wire bus2ip_sync_valid;

  //logic
  
  //Sync from AXI to module's freq
	small_async_fifo
   	#(
   	  .DSIZE (C_S_AXI_ADDR_WIDTH+C_S_AXI_DATA_WIDTH+C_S_AXI_DATA_WIDTH/8+1+1),
          .ASIZE (4),
          .ALMOST_FULL_SIZE (14),
           .ALMOST_EMPTY_SIZE (2)
	) bus2ip_async_fifo
        (
         .wdata({Bus2IP_Addr,Bus2IP_CS,Bus2IP_RNW,Bus2IP_Data,Bus2IP_BE}),
         .winc(~bus2ip_fifo_almost_full),
         .wclk(Bus2IP_Clk),

         .rdata({bus2ip_addr_sync,bus2ip_cs_sync,bus2ip_rnw_sync,bus2ip_data_sync,bus2ip_be_sync}),
         .rinc(read_en_bus2ip),
         .rclk(clk),

         .rempty(bus2ip_fifo_empty),
         .r_almost_empty(),
         .wfull(),
         .w_almost_full(bus2ip_fifo_almost_full),
	 .rrst_n(resetn),
         .wrst_n(Bus2IP_Resetn)
         );
	
      assign read_en_bus2ip = ~bus2ip_fifo_empty;
      assign bus2ip_sync_valid = read_en_bus2ip ? 1'b1  : 1'b0;
			 
  //Sync from module's freq to AXI

      wire ip2bus_fifo_wen;
      assign ip2bus_fifo_wen = ~resetn | ip2bus_fifo_almost_full ? 1'b0:
                         	(ip2bus_rdack_sync|ip2bus_wrack_sync|ip2bus_error_sync) ? 1'b1 : 1'b0;
	small_async_fifo
   	#(
   	  .DSIZE (C_S_AXI_DATA_WIDTH+1+1+1),
          .ASIZE (4),
          .ALMOST_FULL_SIZE (14),
          .ALMOST_EMPTY_SIZE (2)
	) ip2bus_async_fifo
        (
         .wdata({ip2bus_data_sync,ip2bus_rdack_sync,ip2bus_wrack_sync,ip2bus_error_sync}),
         .winc (ip2bus_fifo_wen),
         .wclk(clk),

         .rdata({sync_IP2Bus_Data,sync_IP2Bus_RdAck,sync_IP2Bus_WrAck,sync_IP2Bus_Error}),
         .rinc(read_en_ip2bus),
         .rclk(Bus2IP_Clk),

         .rempty(ip2bus_fifo_empty),
         .r_almost_empty(),
         .wfull(),
         .w_almost_full(ip2bus_fifo_almost_full),
	 .rrst_n(Bus2IP_Resetn),
         .wrst_n(resetn)
         );
			
  assign read_en_ip2bus = ~ip2bus_fifo_empty;

  assign ack_event = read_en_ip2bus & (sync_IP2Bus_RdAck | sync_IP2Bus_WrAck | sync_IP2Bus_Error);
 

  always @(posedge Bus2IP_Clk) begin
    ack_event_d  <= #1 ack_event;
    ack_event_d2 <= #1 ack_event_d;
    if (ack_event & ~(ack_event_d | ack_event_d2))
        begin
          IP2Bus_Data        <= #1 sync_IP2Bus_Data;
          IP2Bus_RdAck       <= #1 read_en_ip2bus & sync_IP2Bus_RdAck;
          IP2Bus_WrAck       <= #1 read_en_ip2bus & sync_IP2Bus_WrAck;
          IP2Bus_Error       <= #1 read_en_ip2bus & sync_IP2Bus_Error;
        end
    else
	begin
	  IP2Bus_Data        <= #1 IP2Bus_Data;
          IP2Bus_RdAck       <= #1 1'b0;
          IP2Bus_WrAck       <= #1 1'b0;
          IP2Bus_Error       <= #1 1'b0;
	end
 end

    
 endmodule 

