XlxV64EB    7a24    1a20R�)�<��55ɯ�aJ�҃�0ٗ��Hé��n�]Àz��C����{<�^�%�o��0�{�|nYHF�l���A�8���T��$���y�Y�3x����#��'��@���jX�َ;V"�~p50����N�Z_�OD��lMp�<\�D��'9��k�B̢��و����IN!cwV�$��Ê�S�k<���h ���E?|R�|fe4Oy���ʧ��ͦZMb�S	wG�%���ٓ�6� b&A��4I�n�� =U
�m��Z,$��8��1����!bާ�
E�W]�j�@�@L?���[���tI^��ڞ�x�dS݀$ć�IN�����N�g:�q�?��Pyc�:z��r$ooW�Ex�*Y��i�#4e�`r�c���/���I0���	0]�Vb�
ǟ8Z���K�\��})�w�c9���0u�����omf8I�O����%�(R�ʶ!N�=e�&�C����X�Q+tA�o�X�dkA�f��*�@��2 �<U~�!���m~�W�i7�T�� �A9Ʀ�D���.��_��gl�^w9^W�k-P�v�̵X(�q�U�dK1�k�
px�t`����D�r�l�T��ϡ�᜗��	�V=�8���fo�s{�;�n�q�?l1Z��$ZQ�����o��Y��t���L)�@A��ɜm�X��u�b��w�<K����_�ii�M:8���q��b�Y���K�+��p���Jq�y=.��K$P��赊���C96��7v�?���?��O��VNp�כ�"a1_�xg�ۣ��e��T��4�AY΀�0�Y������Q�D���%�2}3&��.�I_'S�'d�w�yu�����s�%c�	���[���#+��g����܈>}�q[�v�y��c}iUA����Xg�xy���v�4���N��٘��<����d	�x�*~�(n�'�C�^�%�������!�u�OnSWXX
��#���f*#�k����!(��t�y�[���G��P(�+�M��?҅�a�\�7����\�3�p �9$��[Kƅ�)��g���x�(�(�9n)o��x�-|L����6L����	a{�s]Ʉcb��u qa<r�F�h�2v�#K�Րf'$�W��G�b��G(�[�1���r鴵 ����y͡-�w8(N�_���Sޛ^^##�޺8}��#n*W��xh[�qd7!~
�i�����u����J�(x�6����*�Մm��Ɨ:DTB�n��if��F���`�/}H��d�U��d֢�L�����F� ��1��gg�G��y6.,�ut��,+��j��;�B#��Pt~���B��~�*�Ng��޴9r]qL��k(�h�< '�rʭ��|��У:����;E����C����"�rzG_��ҫg���L�R�$��X�� +Jc"m��t^�j��#�n������Hy��#-kf�>O
��T>��ۦ��68Ǯ�@�4G\�\���~N:��U��g�f����S:�aS`^��M��L�^�v�����@Ýz���Yj�2(C贃g��Q����}@�X8=h0F�@�N�;�v�����y5[l���B���~0�k�/a����6�Q�_��Z�.���K�Q�]�+�0�AnC�E�O�<o��(e�zŨ�TV�I��(`Ø���kCழ�>9n@�T���>��~�t�O�ճي���T��$���Lવ��?����aSu�b�تu�|
wxS@YaE\W遷��'P���(��PC��2��zƓy	��'��nD�k�E��,�@�iIʒ��a����4��.�ja舩\��p�0�&_8���1$.M�}�ЋL�7��[���S��1��+���eǨ>Glh��A��1Q)Q�����4��,����Q�p+�EC��騍��N9�8�b�7�$Z�.���H@����m�O�]ɹ�.F����ǈTOs7����zj.qR�
�B��O!��=�\�T�؃;�NBD��ga'%ݠ�0u�k|�W �"#�#M-���ӂ=���ΰ���!n�c�p�j�"�wd\�ݘ�gb�ȋ�年y�GQ���~��;yZ�%<�C��$��JX�&���5Y� hV?�/�*�b<6$ƀ���/g��
�͚¾ꚧ��^�)�.�5W͒��;�E8c��!��u����auM���N <��%v�GE�"���]H���5b[U�xDL_܇�PbH��?��[���h��%�����K��,\�'�ͦ��}-0΀"w_{�7�A������N�$s2
=��H�E)�ḱ�6m����7��/��v}��_��ꔗ�. R�_���E/f�ɻ)Ľ`�Je��n}�X�6���F�8�P.?�U7�ٟA����0���Ό�τ��1&�i�j���DudN�����،j���cі��i����l� b�1^EV�(�m�2_�b��'��Q�h�G\�\�BX�]@W�(x+@o��V_�^dAo���r�w`�
�t&�Z��sω���[��Z��>v�NM�d�Dye���?/��=/X�ȰU&τ��^����]�<8w��fi�{��Vwg�ܥ������� x� :���0���$"s��l����F�:��c!!���c�3>�ݷ x(�vˠ5e��z?��v�[����0%]����1���.���q��?d�|+Hk.�f�L�k��J���-y�]K pT��H���f�>g��8���妧��]����,TƯ1��b:Ԡ�D]��"P�y�5\T�+F��q�BV��9O��4��2�y�L���b˥[��.��/�A]���G�ڷ!6���u���?��2��� ����}Bs�K>�P>n`�ɑ;�6,��d~	�"��4���8���t�C)z�g�z���͆!܏u9�ٞ	o���L����s@�W@)$&#Dn#����RhB_o~H��s��V0+��ӳ�-�=�k���� -�����/�)zC��S����£ ��c��J��ʮDBjЈJM ��{&�M5g�xfIcG\`y�z��ÚWY���ʪ2Rh��$?Nu͹��ы5g���?Ɩ�Y˷�X
��ٙ|;6X���[�i5�O�����,��Y�`���K9��Kf�LM4��9Q0H�����[�e��a��b�q3\*��Z�	F����ۄ�+j��ǎ�dD=()��vy���H��3L���j��n�7�f��4��͙�����;�!�਽q(����� �3��/C����0��UM�p(b�]���ǻ�w@skpm�W?/���G��1��<{�F�Qy�(�fՌ_�Y�w����wI<��$p'�jQ%I�K���o��t���1�{��"� o��d�
�z� z������69�RZ�^�V�r�ӇӚT��&�T܅V��3k��koeגQ}�����C���Wj3��k)Fn�D|����=�͕�8\r�%�W*���9��9�z����?��>l� @ܹ;�O�Y.Ǧ���c�!�"���M���!�liQ�0�,*��Oq_�i����D�Ԛ%��o���@��c��EFӫ�`�1�F��Kʉ�`��<�i�����S��NUO��F/y|�2��ܽ�2)L-r$[�0H��kp��[���x_�P���S�ᑵ2�����2��ߌ=���B�$Z���i��n^|)��H�!m�a�G#9kdoBov��ȅ���Y%��s��Llr��"�0�?H>�F��6dx�sM����*`t����^�������y˩��
O�X�$���T��l��[;bH�8�K�!����*&w�Qr1��&�(���1$%���Fn����rf+���o'�G3k��V�=2�3�щ��5A���C��Z�� ���
��|S;2����na�v�� F$Ά���f�O�b��g�If�m���R��~Q}��S��y��1IMW��d�1K'�GU݉X�j���i
-p�z�*�ݣV�]���A*l3��F�Ew��&� �M���"o�׼'�@c6E̽��2+�80S5���6Ħ;�zm*�W�	�t�-+�=Mh29�p���Q��X��U}�q|읉p��8�$��j�G���D�\+�|㻯j}�|�dŦxN �_e8ෳ?�l�c m�_]� _9X���'�{�heK��B��������zl��<�XԆ����q�KȾ�<���\��P�Z���0��{��t�@޾�+��t��������[��'F�6V��6D*M���OsÓ_-?=���~/g�S�
�|�J�]�`5�:G����+�ǋ%.	�~	�����! +3��`n���m�e��{����ͥ��T+�%�=��1-�Q�uG�i�V[�1{�p%��l}P|�\���P�af�a[-���tD�K*��c͇�	���������dX=����M�����_�����,���I,�y,��k�u�>�qpۼ�����w �����th�9�򬻥�*}[I�_�y�GꅺAQ�ZDo0���s��،�bMKS�������iW
ϰ����}	�b@���Ԃw���+٤�5�X���۹L�..
[W�{]�il�r��y��C���Lvү& d��RU�d*b���^���E��ۣ���"�U�vP�E�̵}�Zк�R�j�\��,}������ H�i���jh@ב�G|gs'�t^�Z;���%\�4>��XqTIÛ%i2�. �K���\h)�k�s�_}�	���'V��Z����ՓD B��� �y'��H�M�>���Ƈ���7�R����h�E���,�C��0�G�������*О.} ����E��OLC3�y9�Y�1��U���r�����\/'Uhì[�z��F��ô���/�j�����y���QSJ�׋a�=M:���]&w�'J9���|����|�3�?����K���%���NP	2E� '�G�B՗�Y�R4+X,	xM��{�=��� g�b�_ժ��uZ�w�_��K��}a�����$c����mRɥ+�m��y��|���t� g�}��Ko��u'T,�=�5n[��T�]�)�>%��.,�[�������ˬ�G�f�D'bD�_d�4�CE+�B�� �D�Q��[y�Z���-�C�@!�(�%�H��R]�B�ozQs��Q�q�E}'8�g�e�֏��X�PQ0f�� E���Pin*�+�/p��O�*9x��r�T�a	m��j`���n�c|V�\�[���uI�}����˞��g�W�$t_?ZM>��d���}�>�$����C�a?�V��/�B���	��t	Ĳ�A�B����r4��8`)݃q^���6��Bp�_�h_�s�_����ڏi�6<Z�>]��.�<�f�EFʶ��а��,w���9\�T�ю�憇��0e�lT���~��	�����v/z�t��؈<zrs�������w8���Ϳ��c�|��O�P�>�X�l���a��莋P��\N,aq� �\�1s(E�I'%��LZ��v��`�+��j=��
C�yI��`%�A4��
|.xD���0���rs�3_	�Ƃ�ŀ��Ax%_"
���5SmRԼJ+5��Ь��Ɂ;��4=:����qW��[��ݾ�7� 
��#�J(�L���۟3��Zϋ��W:b�oo[__;��l?L	5pD^�BW�|+t0{��M�N�I*߁�hM[�^NJҁ���V&��p%�"H�'����-<��O����7<tL��-t>%&V~ߞԣ�h��\�g�k������1%��վh�	U���.��������N�2�;s�b�DÞ9�cL�u��k!��6����_��
�ŔFS!��Է}���Gd�3f�K���#�0�\ڟ�ء&H��� M�G!j����8S<�Y:�'Z�>#�7�P��S%�1�� ������Uy*��.4:D(��f�q�7zȧ���E�	M��BU�tp*F�>Au�3��6ã�!β��jI��s;n��N9��A�p���<��rQPڭ����Y���)֤� E����V��+�G`�ִR� |�FI� ��r�ɕM�u���jbܒ2�a�>��\�t}�{h���}z��`��Y|靸U�@�Hi���Vk�����6�	K��O���hAxr���u�#���j��-U/h|���tW#S'�����	�i����̼�G����N��* ��n�I�([�_�X"��[�(8��L��i@>O�5 �H<+� w�65uX������o���x�#�K�.y>O��\&�i׳� �͡�
�.߽�:��j�i?` {В,�j�Js,�(��+��c�OJl"� �:��Q@\���O�߸_NL�گ��-P<���C�}�S�9dB���L��M ����S!m@��E�m?��<i�z]#e�*7)���P�S�>�5��I^�,& ��\�X���/������A�����&�G/l�=�9V��Z�����n:�VcZ�_e��(T��RAeOjֱ4mOJ=\��]>"���̟J���W��Ue�&=r^b�k������������A���9��¤JQ�|Y�2���|"��