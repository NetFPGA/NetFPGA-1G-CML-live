XlxV64EB    fa00    2fe0] ęB��&\d�O�hަ��I0��$�%����N��#Ӷع��7*A�^���#�>���;�<zƅ'6>��A�k<��F1�68�v�ӓ�u'���2E���FB~�=��7��2[ UN�m����q��`�z�<���>-ki�8�s%z"fwsh`&�*�c2��n�_�K�	*g`����jMCpܞ(�GRZ�]Lii@V�ľ~F:g��hj��֒,ᷤ���� (�т�� w��Ft�6�#(�x�M`$oiݿ�2�̆� ��$�s���7����Țy��6܊`�T��_�7%�p�Ň���O�S�����O�R��=�_��x�"uu���hKS�"qC�5�C��E\ǐ�5��2T��%�w�N��Y/���F~h��5X��
��h���F2�c/3���3�ڦe�,�o�s�LX�f�4^�<�Z7h�߼�I}	T}���2��`$�i�˲���s�;:�9� + S5��U�l�nX��o���[��� E;tu�l���k1���ͩO��"�`F��c����8��V��&�q���u���
��*������ᇴ�F��h ��4��� ^�w��ї��Gma��]�9��x^Dn`���yb��F�x�P�Xw������N�|��+bIB=����}�oQ��KmA���햣z�RT�o.}5���_�֪�ɻ�K�G�K�5�>-�ĽlwPw!����CQH.D}"�ɞ�y2+�D���o�Hb�U]r
��z*OL����W���L	����9�u�9��	�η�\�I`�" z@�/|9�~�e��b뜁a���:"��g�1������yl�'�ܼ�̫E�gds���:��]��"��0����A�K�qB��x��L!L4��Q�V%��x�<n���bg���`��B�(5u}��Gv�3C�G�������67$>���0��F�Y�|Fu���}��9:���"�LeR����0P �1�Kڃ+-0󌟫)�`���	�U�h�`�����} ���r��AI5h�<��9U1(�i��,k�J�YM�V�ۊ�L��� +�!e�me���G�V��Vj"g�v�;ߡ�f#��/=p3!ZC�� �B�d᯷t��G������a����ѝ��6�A"�*���?{�}\��{_�G��}�
�X�ⱦQ�泪P"���:�<|�������,��i\ui��j�a�GS��b����n��=��>i���P�yJ懳�-����Cy>�ȩ�1{�d��%9��ه��
b�(h7��>�9?�6i���&jƃ�.$���h���s
dN���"�%+��چ7"'�5�l�9fpj@��Ҕ�\����n����/B}��V~;����C����o�!��!'4q���6��m���D;_2�s۽����5d��EA�d$
�z��)�4	���Vt��8�*K_����{��!��I�Jߓ�cx;�FCO}v�x�t��,r�-]���d�WlΖ�C %.{��.n��Cbk�}����a#��7k�uU
�G����DVa���O(�8V���FLo��*�x�-����0,��~�Im�% t9��Wwd�u�M��=�L�`�t�S7��X?91;�K<��ɉ�l�?�ι��}9����y��o����)�o/#��5���� >��V�''�9
y�>ϴ�KZ�� ������H�'�{l����%��C���-Qu�Nc���ҳX[�=/~L"�J���/����	k�~� �y�q�}�LYi_+9���7�r~0;]j1�KWS�^Ū*_��o�W�[��Ny�c�ۍ��	<@�
�
.�"#��_���o��^���r��1�����F�
sb�o��{1��?vE��A��r%��P&f��)�����iWq�q*%�B/��o[�)Y&'��'F�Z�Rg���,��@F�;J��Q��Ρ� �A% ����� ίH�Џ� ��:��_{-L��'\�<5 Q4��v����R2���Iڐ��nW4�P�+|>�K�f�-�E��(�����5&"(�9bx9�yEq$W��l�����4l+b�|rN�sڼ.<�<WS"|���}���r�h��>M�Lc;�	B������3\���� ����	�4�V�>0Y��h���IR�?��X�A��Y��X�?��'^�병�.|I�e���";��`Ң�'���A�|t������*�ԧBG\����Õm�}��<���!=>�Ae�y4�.�C�0�|	��ߔA�PҗwrG��"դ�?�.r���#��9���;�ǹF����=��J���T�S�Rn9��mh�X�v��1��kx+����J����>�Őď��ɢ�I���ht�:��SQ�}OƾCSs�l��c?�B��Qz��My�I9��_�P�p2�b����G~�sW�����C>���ibPaᑢ����.0Zٗ��P��h�1�K<��y:�2�d�7�9�
A�+S��t�ꋇ�SYw��Zʵ�d!*wć���&��w���</�ӥ}B�B,��1�{��SM�KNRH��)���G;e`9��Vw{Ki&��cT�0>��H��[�V;8�ښ�75�������ܸ�k�=���ŗ�<|� LV�)��)��N�+���&�$��u)�a��,���@�@_��1u9f��̾�P��m��q�!$g�ײMŏ���ܵ�6����������>;�-;�i�`�8"44zL7�a?�T"�H�3�JX��>$e���x����\v-�r���_1/�jaU$����g�*y�0�݃ݗ�B��7vΆ��(p�V��8�C�J�c���i�W���g\NX�FSN�q�H�������X�_΅bu�?7��o}�<��R�(���@a�ƌ�=D�$W>����{��D���u��X�+��	�8H�|ل���"����?kS�u����"�z��Va_�`7jwH#q�L��F#.Kɴ�S�f���P�y�s^	��i[p����Q��z���p-n��H�_��|L�N��ZF52	�{��>'c	"���"�:-'��K)�L*tQa3LX�5�
�!-lL%5��L=��P�ߖ�W��mB�N�.;���	`�f��~Q��;��`�����i���c�^�dl��y@�n�h�SW�Xi���jۧ:�Թ�İ#G�g��3(��J���;�b������ߴ���Rxu��*^֥B�����D-��eP�yD�&�9��\1N�E�=�3�ߣN� ��+�B�I��RG�̙rJ�������pwmB�c�$����K_���_�Fw�Kh� ���D�Ÿh�l�j���h�@ju���60��H����1�zK��9���3GK� �"�i�q�h�����Z�P�{�%���+�����Z�[�YR�l�-}ץ��(p����^-3pO\��m�$rz��"�Qf�{�>�KηUؠϾ����Ղ�`]��,VV'-3�:��D��@&�L�Z��fj}���Zo��������(�,oB]��w��'m%@S�t� ��1� 15��u_;q;����7G��wr+C`(X������!NI��l��Cl*�)f)VB�}�)�2��Yô;
!@��jOI��A��Q��:�UE���z�t�yv���Jyw���:�0/��w��3^��q�'x���.s�j���P�<�X?�����r9�cYd3~�i�K�&)��YI��������>�˵��)�F>O��v���mV�q����0u��)[����e����P�Ͱ��e�f����ȳgWaW�N��%���dQޡq����V��<H?�j#�'ɝ�"1�ŲO(�"<��3n�C?w.3\��{��/�
z����"��
�ޥe5�o(�D7�C&y�ᘀAhz
 �~�Rq�*xz���"ޠ�7Ϳ4���$���t4b%.`f�����X�^�[Mfn��K5^�v�BXl��ɒ�f{�!C�G>Si��]ќLI�c���ߘܰ���(�q\�[��4� ����?]w�Τ\��J��&p�g�=w�6�NQ���}��"QP�v��Ԁ K�h��h�L���+j�R!�)ѽV|yv��(�����iݼ=O��/�PC[�_�=<�p�*Dv��=��@k���|�J�� J�7� Q�U�sSc޶�c"���*���BK�T�Q�˖M�X5��VT�ҁ/	�.ۮ�j��~Y�6ƛ�ɹ��H�K]�OL�"Wfi?� L+h��Q1�=���E���/<�AV�qٝ�D�嬁���nG�g�^�4ދ̒���܏Ƕo�$�q�� �gT�A��!�O-"��ȍȉ�Ԭz�A��-��Vf�	H�)���Y�p���Ӫ���&���*S��uAl�Eo��+�fI��ѩ���b��ߓįUPop�^��"n�s�`������l�b��Z*]�V��
 B�bs
�O����Y��E�\��t(YG�PZ�4�2q&�Y�+	�x�@.�L��7��B
��A�O�W��V���Fu@Z��,��pбy�N��!�s�#�-�Oi��PS��,ޚ���`�"���af��g�BE�l�}L���Q^���ֿ؞g'آ���z%	3	�W/����t0t=��g0�zl�`戓&��V�a�D�#�����ο�$.Z��:�V�\;��XH|y�j9	И�;�w�˷�=�Qn.�&��T�b���9jy# �i�ҵG�mKCEH@t����k���v�}=���6"W�( 3V�΢x旅%�W���� 	�
�ƱwB��'�䳱�8���H�n����I$Aڋ����|w�>f�v�#�A�	�A�0�[���I��~��������U�,\?&U7-Us�7gk�x���5m�ŝ�Ҥ>!9Hr����[YƪO(�AP�sgȈ��,�<�3ʔ��CF����i3�*��S�~A;�%���uMA�!\�z3[_b��iHi�v(�v+�J�=���V\3=+����;��r�(^1VաqFqG�\r��^;"��څ|��\J�s�@��,$?�g
�����Am[�,U�� m6��-�c�y���e���4�sf�Y}�h�ڞe��W>^LLQg�8��r�n�?��y��6"\6�}_��6�-��K"��S��W����3�������V���f�/*������rE�
�	���F/���Y���n��:{��p�NX��d^�����{ҽ���-��Z�Y�K�AƤ.sW�:A>��&_"��袱�G��#6ܘ�@y2���� ��gS_&DZڙ錬j�dզ2Y��O�fxl�O|ݎL 8�/Q�䞗��kZ�b�mW%��ɵu~�[�(��4��\������@ ��%H�4St������?�4��N��qw��S��Fc?�= '4O��}�6XT���:���O��<Q�ʬ���2U����fs���]�lJ�7�>��Ql���v�v��'b���N��vK����n�Cv���������ʜ[�poڰ�W�a��?����g�|1�
y)$	�%vY�ܑ�L�ت�t9���'��]�����s�R�Q���/ ϯq�q3W��MeO�|�c���\CX����m�j0�����C����u� �;�D�V#����϶�����^������?��&�o����{�1�#��x(dև���#���l��r���.A��w�y?gS�� Q�-��$�R�R�OFU�I���"쩋��HoB��Q��}#�;�W���v��k��/��l�$��@�>I�[?y�cu��s�&��g����"Є�U��� Dc;���Ml>l����5�F�����p,�nq h^�������2^�fV8��ї̾הN��z��Pa_�,�Η�&�|���-U�3��(�V5�i
��>Y���J�§��=�_֠���C�!U;.t�BC�q��Q�m�����+Dw��z�6���aF{��8���:�&G�	���@F��j���K��]�=������Ù1�P̙�<��f	_���.�U]�]u?=�)�\
�@����q�����	3jv�,`�ľ��C$╆��s�/=�\��ۉ���n�	A�+�Nǚq8�M�v&1�L2\�{�������=17d��j59d���_J�blaW���b�GU�!\�d��(N����B�?�"�{������"0��O�ciWĽ�F�*s3��̄�"�A��.D�i3��O�ZL!�l�J]Q�����+�����y:���a���<) A㳯�Nv2CI'qi���Ոi.(��7*}f�-D�+��q���X��`�[�,��'r��P-BxynhX%	GU�`���MR��g8ҡx�c��R��0��})����?�O(Y��7�;+W����C��=6��_�4<9
لR��z���7s��I;��ޅ��m��n�G�[��!}�Fh>� c�g�[؇�_�z�������Ź��Dj�Q�~@�M�L�T�T1���n���ID�`�~��W�ŋw0�ʕf;~7�.r��h]er�K�Z��B��G˹��u���ݴ:��${E6�������"����� f�|����͕ C��L�q�+����f��9pj	{��B�%���O��3I�K@�жRh1�
��3mei᷌3�����Z����������`P�����0�>�M�Cok�ĺ�����G)���E��.�B2%����g�S���nU'���'�jL��[b�nt�ϰ�O�NB��b���-���|��6,��qٹ���P&�J1  �3�����v,�����+ y�z^ ������a��֍�+��p� �	����������'2�&�&�y��2�(ۅ�I�|�5Ł�\��+7io�[%���.fN����"p��Y�����1�o_�E�����v����^�x�0]�����Nopt�W�����1����:Ed>�p���'�O�1kid<�{H�Ύy]�9-����_}�|~��Q������0浒�f�������o��/����-D���!JW_#_.��^��z��O�o>˷\-�j&-l�<�8�I�V<mx#�'.�.��ǰQ��\yMYT��\����>���ߊ��U@���t�a�|X� �q��g_9�O<~��9Q8_���^~g%~}f��\�� ���OR���������)��)_�9#qx~�^D)�80��۟�-e��:L����۰�8��J9��Fl�w�'fƴnv���P'ޔ�u6�X{�;qR�)��5�OCt�2���_F�)��XiӽPeR�Ϭn�B�+�I-\.��e��q�-�Fݜ��Zm%L�����:"����æ����A<lR�D?��yLe,�	?�y�����"'Uu��u�'eg���r�	��b��-\Ng -$�~f��ࢗ�$"�Z���غN�;a�*O�)D��Y��X5�?P2ڛqS~&m�X���(3/��؈#]��܆�>��.T����!.��Ձ O�S���)%C�%Qf���_���&R�U��X�����6n�+� �0)��ZJ��w�m%�r֭��-����'R �P�k�j߹��j8tī�GP���v��҈�g��=	��f|>Cn�~r��R��Q��+�M+zx�� ��y(C0I%�k��l6$�*�ʯ"��4f��]UI��5�V�x^^q)�ܚ���+��<���>�N��ܒ^ܡ�>��k PВFr��	h�_"��q��,��<#�w+ �A�}c��\`��� �u�?طr馔/�*��!��/k?U_��NBVG*~�+�9�{l�4��B���撣I�<G��i/wU���yVHZ��~��0��h����a��F9Jx�9�|��*��Z��u�hsv�1QvXve���|������x2�o�M!Z��UG���a�c��o����X�x]о��%�F8�j������%�,/��
�8�6R�ȟ��ܭ�U�c�2%.�xt��^y)�/�h>=�h���*�s�[/*�W.G%�{�D����k������Z�D5kB� �_�4�]�Vnp��k����������D$��:5PZ%�;�r{� ��:b��'qVt�6�6��|"���po�B��RoY� y�����DWJW��㐀y�d�b����[p�'E�x�Y�A^-�ϝ 6��]���yi��}�9ݩ����}���=)N�|Ҩ@*�������H7|�:b�d=�~ǉ�$p�c���Q��5W�M@[��*�L���Te�$n��Y/�����������mA�￥�y�vz�s���G�����F�O#s�C7=�x}(�6{g�j���"���k��1I���N{O̬�w����j��)�|��ޤ%W���w�L�7�#��5,�5�Ϣ6�����i.#���kv�j�#�F�2iˤǐ~[��H-��>$	�wzQ�=��iMyy��\��Me�,�5fD�Ev��[h�x쒨OA���Bb��IV�r��"N���dL>�n����Dۺ�"0��Gs�0�����!V�/��>|��c�eŶ	Լ|���s��3�֚m��D+�%�dXD��'2
%�><�F�=V�/|Q_F����8@��f�o�SR��~!�O�E`���Khh����%1�E��h�K�5~��ی=7X'���P���t	���ӯ(�L���/���JJ{�Z��b���E���lu��⧌��[ƘV���N�5ח��E�&��`�K�8���R��v��5��C��lxyt�����Ffu��E��5y��C(y� /1�`�MWN����C�C:V}���rB�RD���a2l�#A��`BR�?���͠�?�D�Mz.w��s������`D��'��E��{�ؐ�"�?#�0ב��B�rX^e���]``4��/K���� }�Wڳ���ȼ��� P$���փ�Iʂ�����
���(��� �����Z�Mz����$�����ls��o>�����M��!�I�p���>�����s�(��-\��!������l����AXe	�ە��̿j�4S��5�{L�9ef>��ss`�b1�˫-p�:O�5y��uj�!
o��*��q��	��=��#��=0�;O:���
P�Z�vvY�"���J�#d}�ؐ%3�'=ԙ�X4\}h���������)3 �cqH�2a*�.�*���7�F�m���vq�4P�e;��;���n��ū�����
�`xN�	PD����w�/���مS�nP\����ڱ�7�ž^[��/���"�[�櫰0\}�̡S�~��V�� $��������8 	@�3$������v	��."���'��0�R�u��#\��em���e+�vlS�4�~�/�C10�U���%C�q'B�d����/]^����d�8���7�;W��F4'N_#��Z�3iφK������7\>}��s3.���]f�����93먟_�1�Rf$��mJvɆ�v������>�slVRd��$sr��ᄛ���Z��ڗ��,�Q�N�AW {?�Q��0�����7��bpc�
z�2�j��p��YMa&oBEc[Ur�6����b���l9y!�^�����>�L��ٛ�f��#ejGT��B��<���5���y�06]�=w��bK�_��J��q#�����tw�ϑ��)��Riɨ)CV�ɦ̠_2g�(� �7�EI���t�M��o�P���T¶�ѴZ7���%3m��ឣ˚_ ��+��^����\a�D����ը�t4zT80��Ř%����*�5bL��UP�)�-�7�3� j.�Qf�>�G�����>M�OvA���:uK�� �dSSj�y���8!�<��1�5����7Y�?g'nq;.���0�t_~�n�N�{��ϣ��ď��㾆}W�t$y$9#�e�-����j9�&˨*�*�r�hM��w��d�'-��	Tl��Hɏ1���F��[�Qj�\s�-)P�-08��k��\sG6 �Hj<5\�����E!yN�#4ǘ�0o�/���Gc��Q���$�d4��i7~k]���sצ�5(����}�ݨO��ocF������:�;�s�Ȇ��� �s�~�\�NM���H����{�>��������<���<�z�%3�|�k�$TR�E�ԓ��0��@���k:Uh�D��Cs�ŖEgtēB���on��u� �g:�v3N*�kh�рY҄��d��R��=�DX��'Y�H|+�tsm�M<��	h���C��Z/e�� �����ׅ�o�QKז�����lM�RQF��Ǫ�\�A�t�Щ�u���ɂĒ���J�y���CM��D��Z6K���s)Zp��q��*����hTSE)����쑄�j�ϝ�g��jUD���#
�_ʒ-��Rict�$�3��Nn��tfJ�Β�� ��ve�誠�N3|�F�����P��j��Y�S�n�`�?�Z=\q U�azZ0�)�P��[�^�;"ҟ �g8�>�	�{�f�Dv�F�Z�uc��[������ƚ��>���,�-�H�������z�ݝ��k2��>&���~P�b@(J��V��|Pp��`��S$	��I�j���!B����m�@�|�	�0�Z-9kM
�Y|��b��׽�Fa�3���_�:���(Ѱ9���B�@o`��c��ܜ	�Y��4�:���0�I&FM�lip�+t��M���i��o9Y	M)���qwV9#�ΫG�v�W�}�8���R�l��	 FK�K�e��eҁ�K�x��F+�]/lpV}��󨔢�g-_��3D6�ݞz��>���94�o�����f��K��e��ѝm3�vf�e���E�1M(yH�����&��vGg�
 nֵ���_jQ! �e���q�aә>�%�W�>Dիf�Mq���x��I;ݿ-L"g<�k
\D剌�n��s��$��WeZ���(~ų��GŨ�3�u��MVx��I6�a*��حW?������`OOĳ�Ә?!���,�c6�����b�1kt Z����"������M]��k� ,�}� @Y�mS�Ff`������6Pq�-O,��t	�6��%Q"]O���ٵֺ��~�0T��`؜����o.�����n�[Ovd�ny������W�(���ڬ��="Ϲ`H�F}�^�d$�4�ڗp�2(%��UK�f{'6:�;�b��ǋ'�b�����|��'Ў�i��ʽ=9
0〩yrJ콫8���u��ǃJ27*s��7/�8*I��C�5��n��z�v�:^q �9���[��gwmC@��n �v���ܐ�L�.�m"�F���4t�+�JZ��J���Iq�����U������<�!��hs�3���h��)��w�N�
a��d�� *\���.����kC��6�5Ŷ�]`�/h�XXS� d�Ta}���y)�AU���BRʋ&�W}8����&��0�-+�6�vu�D42����\!�H~TW�� �4�J ��41�0k((w�G�ʺ M�c+[� /��ŭ,@�(+����V6��� Ż"ګ:���ι���~� �@m0~�y����6:��e3g��Mw乛�9o}ɥBL=}Փ*�g�㟟�����)�L��^$(FE���K��_3�Is_.��
|V��u�k`�?YR[�YP
��M���W.�n�rB�7߶��	+��mI
���N���L�C!xD>j���%z�<m���6�V�n�Xm�>Z�� Z ���/�چ�DZ���*��9n����"O�Y.�Ȟ{c�T��.x�`|W��������Y��	�J�^��hC��.�a����Q'�-٦�D��2~�X7��;�!��{��Um��λ�V���,$��S��
����U���rMG���7���,4o��R�R=S�H� ��w� �wl*��H��-g?����:j�� &����8��ʽ��.Edy=���.N�v�ͳɫ��G�%��3���-�It
����l��� �{D�Z�@�XlxV64EB    5f88    1450��4#��-�a	�u�{��?l�vG��G�����(����K����PᇸFƉ=�@��Γ�N|
Fcf��n'��<��Fe��������]��(���G��L1��&f��L��ף�Éw)��MQ������K��	�'g����.�}�S�3���?�e��B���>G	�!#��Ɔ<7�D�*�-��6R ̋H[�Q�7Q���@͟%'��E�s�2w��#-/��0+��T�y8p2���O�GS����ׁ���	��� �76�ʈ����a{�����xAY����g�'@+����ԀE�Y�Wr([���;Ӑ6�"��v���Xs�mGt����
l����šrZJ��cΧ{�7�Ȣ�1oMݨ-[�]Eӽ 
�U��=���Ϟ%�}���n�[x���mY4ih�r����<���Z�_����o��1͆�{(#3	eF���gi�O*�X����1{�)f5�!��ta�)!4��*�/���˴�V��2��f2js`Ǖ��E4=Vʤ��L�0`}?aUg��3W��=��b�_��(.Ad�v`�̖����Yi�k>�!���#����}��}S@��כ�o0=c,��*$ܖhh�� ���O��ۻ����*�d4�����[�U��_�dO�wF��WI|]��ʇ�G��D��]RPhv�S��N�*��\�W� #t7�VP����ff�ÊեF\��xԞw��`��w?`�M��D2D�ԑg����g�x5�
�[_�,�W�pH��q��P0�!�ְf�8��i�㫀WK�?$��������Řl����?a:p�E_6F��8�[pO�/HH6J��.
Р�O��6C;�v��p=,�tV{�K&Ao�|�p2�A�B��g�
e=�(�s<��M{��Ǐd�p�P-se�i�<�ݢ��S-nKPìq�'S����Jڠ�kϬD�bK�ڀ�#(ѹ֌�h�>��e�a{�ӱc����5���-u���a���}�,��׈���I��<�|�:��I=s��xwPtQ�ʘ�@~,���s��R��]q7�â�]�'���񯒡���}�7�_�I��bd\G���tn_s���9]C�Ӥ�Jf��!c#:�B��7)n����^j�GQ�l��
zo���+���yc�UQ�%��3����Ax'��Ը>���z(�Em����X?	�'�`ι�K&�����υd0p.�U��19,�N#�KP�"O��cc['
�Â��+�����:�֬Q�(�����V=ϱ����.�����ε��IT�L�?���6���̣�� D��)ډg�=E�g�l։l@�3��zdfA�)f��ni���JĐd�=�WydM����!4�(�q���*|�V�G�Ĩ�q]��
�&1VY�P���R��d�� |��2����O,yn��݈�D��
6��.6Tc	�8���Tw��b�Q*��-����<ɔ
l��,g��Sܬ����5a����Vn�.t|-^�<Z���P[�0��i�(7���&�*r�� �=�U �+@���pO������4� -*)cg�ѓg���:�qG�^��83��/���>|���
��MĠ��Z��lW���x*n����K[�~��Ɛ<�c5���m�~S��t.Tm�*ͨ�:�n#%�3� '��_��%�����)(s�7m��~���^�o���*jZ��
�@�>���[D��a�h�����B��	X?t�'Jh��������8�+������ZD�9�2r3�YL���'a?ɹ������{�����n~(��'FQ������byv�M��#�٧!��K�.��>AD��;-�����h�SM�Cd
���r	��	�y��0K@������P�X�^�cP+��^Љ�������3�db����:�0�u<������9����q����X�f@��eip���YJ;�|�C��k��O03,�^ja�6�:�	e�����ax��\��tq�_h(�"mmŎ�v�����n0n���'!���EZ�����#e����{7���YˢsK{t���U��� u�*r���E26_˂��]�����������u�Ŕ�2��.�%g���G�����1����U���V��m8�
ְO�e�!�S��G<ߤ�Xӝ䌁�2�Ra�ӽ3S!���+#�<�� �w���d�!��;����v���S��m��j��vmr��.ܔ�����'�~���[}Iu�[v��,��o�p���:�F��`;�AC�D��bi�fkl�x�:�U�K����8GH����c6��#��*T�oSpaA��*WBq�5_�Xx�"�D��m�ez��,�p�E� I%�� �e�� ^G>�cZ�+d���|�SjPk�7���e�q㥚�_I�v<ڂ�V�x߄��M����>���p8��yu��vz�55:P0W��p4�,��#t����K�hZZx��Iɽ�2S��EU�ϼ��7���'��l]��ʨ��V^4{F�:�mAN�V�U��Q�ѱ(�қ
u�(c�9�� 9��l�K���RA@0c�S�YBr�L�;J)o��9<D4.t����:/��[�V%&pE� �z�:5m��Y��IF1<6�)]_l�J@W�0j���1��I!W�����Ě��֮���C�����f�7�Y:�1�z^v���᯶Ԁp<T;�G�<7�tf�����(s�|���z�ϼ��q@C�Q�Xk7S���Fq�Z�%/ɐi�qF�ŷ3Y�x�-�tz�t,����5�A|ÄЇIѺe�F���g0.��%C�=������&���@�>�F%���l1�G��a��-�$����aU���R�`o�ңz�ll��X��Y�������v{G���y�!�/1ޢ_T�ì�t?3T�5��l��\�UX�v���}�$�T��h`���)����90#�_1���[x�Wn��J,[�)���*_�ڶ��&#�!�n���p��G�ÉA�@	���"��*�=��Z���z�t/�����&]YXs}�v��O�1�!��z)eՐ[]ElD�# J';4�a\9����|��z�jP�'2�Vv���]
kQ�h0��d.�P���^���~�{v��,�t��9~ET>�N,�,T�L��.���-�R;��ɜZM��1l�l�%�nM�k��5v��9����_pl�P��:�Q�ƨM����=���QңM�Ii��^��.��Sm�����}#1y�#�"e�2
�&V$\��+;�`艇²��s�S{a��tUF�p�i����c͗�O�$dU�'퉁L�`F^��o<����6-���zx�����Q^ȂZ*p�!�������V���%�b�&�j`Ecгm(���lZ�~v ��Sϭ��{>�2/R���H�S�"� ����0��̽��B�T)�^�>D��������5�g,r)e�g`	Ă���7:��w�up�@�Q:$��u����\�^Q�Gų�c$�_�^���+�<v�h��R�5Q��6&�x�ʙ�?.���u��ae�6s���(��	(��+�%�P��v��H���R������|���0�<l:U˪���0��)�0;����1��"�%��<s��q����Ihd��}�a�b��x�M�p�� �"nT���D\��Ċ-}��2��fJ*�P}��$����~499�=�L:��T$=G�B�5�f��J���8[�^ ~麑�%2��l��R�i��usnp�M�	h(�"qЊ��#�*Q�\��HĬ1�>�!CŭF�W���]��A��t	'����N^$���!n�'�tP#r�:5mE��j߅���|����'��jH�0�����^��p���asơ�՛|�Y���x�Z�B⓰�)߿#��-Ax x���)�_՛���� #�{)�i��>U���S��jv���3�脺(�'w]m�x�P\�@kq�Q����e �+��-�ZG1��k�s�#$��劆�����z?x&p�Bg���f���,����](�R� Sӯ�g���Q�Ѐ�{r���W�_T����8��|@����[_JZ�`����@���O��_��[d|��@{+� |�Y$���+S�j��`�'�u��i�bƸ6x�]j�N�Ƨ<�ɟ���4x�Һ�하�p�Y��vB�i�?i�0f�A��j�������c��	�yN�pZj����|RA��5��ێ�>�up�mo��9�?p0���x���*��x,�&�ݤH&>��h����ƨ'�߰������p$�F䘗!�-q\��lLˊx�Z��/L�S��˖��d����yz�Qb�z�g���XU���v�L�������;ſ��e�2�(VX�+��D��$��2�j{�'��C�6S�4���P���R�>JU�IO�6�)�W��M>� ����x��.┑�)��>t2`�U��y���p��j漆�%,��պ(f{������H�XbhI��ŧ��G��Qt�?�P�m��gb>z6]١<���d[�I������Wmȡ m�u��C�O��< �\�a�"��w�)Pr���f��xa����#���3)Ɖ�avx⏤�r>����s���ߌп����~��7K�[@�X$+�퀳�4��R�-����u����=Ի'O*LD)�N'J��s��A^�uT&��=�5b��=~Y)�p�޽�\��f��|������A@��=���F��(��Ƞb�e m��6ٹ�[8oM���9.r�U<�S�l�B��L7����åˁ�I�)�z�"c��  �}���ҕ΋�G'�3����~(��53yA�����Ǫ�9���IP��u����������qr���4q�ǤA;�6�|l��9�,ۼ�>��ܭ��F�Ow)V(��#ؖ����me2/�*n�~�Ƌ���	��}ۂ�r���HAo��P$���ܛS̷?���S��%��Q���nV���<�W�'���8k���	��h3p^z"�`.d��������;O� >s��E�!��,o����F_����~�uL"�d�|>DqM��T���Ud)���C�iƨ� �