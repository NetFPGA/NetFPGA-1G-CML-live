XlxV64EB    1e16     a00(��]�ֱ���X�ܵ9ќC-by��@w�6  ��S��+]t��u�<Aq���b�!��J'��s����g�+�-W�k�p����X�x�<���}��߱^^*xrv��,�N�q���<���/.�܊�X�*��2�|��XW���\64I�A������fJ�c���R���5�K;�]�I �'�B�Jm��E]{�TC$�#���G��r���D���)Qn��ž��k�lX������ Z�4�@���mJ�f����K�$�N�˛��%�K�i��_�����8���Jv�2;�0��+�.��=��(�Q���焸�F�T����;ҏ����?� b�� aʭ����y�2b�f/ra=�t~�[��S3�����?-��bE�ٍ�XE��U'�D[>	�Ɠ�cN9�"�������"��.��_K�����ؽd�Tb4���Q7�#߇iLd��:Q������I+1�h�2�s��!�,IF0����:�pM��.��qv�)�+�c'Cڧ*��V��� d��1N��Abѯ�M��>����
h�zq�pfP�\)cJ��'�����5������l�cџ�6�U�͍�c�C��Q>�>�u�<��b�*%b�P9ŗy�l� W.���TC���3�-T��ZL�Y0T.}¯���L�Hl�饞�A>�c�N���ԙ�E�����(��hJ�Q�_�Pzh������
�Eb�#1~�5苼�/*h%�i %��41p��oz�ۺ�`�k�!�_Gz��
,)��Ơ��+f,��������Ԧ3�XvN.-j��BwD�d�U��c0��\2�S��>��gT�T]0`�/���|B�d;$�ND�aG�A|�eōC��;af�UM���1����@[�R=�hn'�ةV��$1�GQ܏���BHb	�6X��t3w���iJV�%*k�سLq�7�J*��Nb�B���u�ڪd���XH�҂��A."y���">*.l��)	��uh"�V0j����Ei��S��<� I(!*����=(��V��ũ�zr��Qh����!̀���)�������DF7��y*J�#�|%�Г�#�p���u �M�A��UXH_V��ӥ�TK/������g�'f8*����@9/�1�)�*p���DI�@��9^� ���qU�,��� X5TY�;����y�Qр��@�H�g�A��W��h3�(��_W�',E ��)�!�3HY��( �y�!���MԇW)�6�,�4A�=E��-�{i�V�F1;7VFy��US"q�4+Y�wݛ���]��p�M���'o�5q�$�˃�̿Pő�y��v�����}鷥�������^w�	�N޻$P�wb�"��D2O�����W`�H�ޭZWȕ M�=$�dj.v��$�k��lClU5�&�x���S`��e*>� ���R� 
E��+�3ЪDj�e�vW��ߡ⮵��Ar�_\B^�p�"4�]kB��@�KP/ـ!�@{)&�T#Qk�;-�钾�s
�qb�#+���� [lC��ֹ�ml�[=0����"-�;�uN�}iC�s𨣺ˊ�rz5�5�2	������R�GI%�@�/�biG�m���(3b�ΎkD��IU�Yڌx
��=1� ��!cMU�2�p�!~ز�~��$Ƙ�:oTj�b��~����沯 lQ��jED��r��l77�?;&$ ����7=��@��e��D�&e�ĵ&�w�-���E��E���L{��T�ngE�K�<cq����Ѓ��'\ǂs[�c'�'kѮ��"�a����\=�a�*K�A.Ċ�%�<��>Mz�����W�!�q���0�R}a�BHrZ��) �n�\Tj�y��k���#���!����c 
��3�q:�������(��N�vX�F
�p�N@�{��hs"}\wv�i}!0�d���W��U7S����T������q�rc��pFc����0ɝ>���0��mO��ܗ0&�X��7c�=��
�GK��?�KK�KL0����*�_�4��x���%SFB�� S��P��n��C�JU�Ky�6�q�i����ML�=D��!���6��/d�p�)
�9��0?j���5hI+��8,�U=�t�R��O�2��y%��O]�m��w����WK�@~���$]����'���4Vޤ:�TA�^jƖȖ,+��^���&S�~L��$�iuO��{�޶���E<.X;���1��{��)�Q��\�K�o�V�B�X�M�&>�2���  4��i C��J$��dfc�y�ҴtU�BC~�a�l�{�t��w�[;dL��B�X���N��ן�L5�_��X1�J��ʋd�Rbv`8o�ٳJ�§�������I�0C�
����8�:����odI��YD����3���� `�����SI��O\oet�V�xD�����Ѐ*Z�`l
L�6�!�ꊳN8Ga��^#������=�y��>�Vc ���7�()