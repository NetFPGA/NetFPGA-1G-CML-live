XlxV64EB    58b7    1210�����*GE~S7�[nҬ#cZ�̫���������?Y�"K*�������M�'S׿���N���H���R��81n�И�����hw�S�VjV��P@���c��ȋ������l�:�t��h��;�i�U��P�pK� �߭���?�` ��#�Y���CQB����(̀G����alh�U�h͘d\�}�꼟��&�m;/�nw��J:��N�S��\3�0a,L����Vm!�>B�`��(�
z�Q�B>���6+�/p�Ĕ�U�Yc��"}f9�w,Q9�>�� �����`Es5tAp��s��7�6j6�
��v@ΫX�3��*d'h{��%���-�z�3��a�� 68�K��`#�D+���Zj�PwjV���r��\�ޅ��YHs�F-���^����d����� �E�s���P+mcb3w���ф�ި�L��H_���]	˄���h8�U���໤�\���$WMz�<GH���og�[cS]���Lm�1$[K���d���i����(�� v}�������z���[���ȏ��а��ȳ��u�p�?��m��ۚ)`P"<��M����}ę���j��o;���Vs<rz~���2H� �����˲���i%��LBb���F��Ћ��Ɂ��c�1�Fz�+�Q�����n�q���X?渊U���5�L��rE�43{��ϼ�[�?��+G�s�(�P#�cS! 5Ŧ�e�^OY+}�<؂���!�=F4���8�%/��"V-lv��X�[�NJ,�����z@�&���웭��/�������#d��R�E&yn�7{r���rC���0�䊏	f��ʂ�D'��USD��M�f�4;i�r�x��o%P�q�3j�-mU�m���_$�O;!� M�{D���-g`�z4* �'{H�]ZD�8�u��?u$��*���im|z~�nDL�����{�'Te�GI�}��M��� ��9 .G�Z����"���Cg?��*k$V��"t�5����y����t,�Ty�bc0�VJ�j3�0I���%v�G��Y��R{��r`�0�i�
27ӱFԍC�lU:�*���/L��8IC�P�9-��Hvg�~t*��iH)�IIO~�&(�_��Rc�л�| ��@_J�8�����֖t-��������Z6�U�s�qg�VS�W�(eG8��q����������l�=�l�]̾�v�'z�Ӹk�F�6Ai�f�/*>8HN����|�_Kb���Z�[h@���f{���g�a�Α4��(�~&�!��������KL:I�9N���J���f��;e�oy���SD�4�C~�� �EkK��F�wܛv�Г��7b��M'm��Hpn���j:��'\A��M�,1=>��a��%�Q��{��V1u�{}���X�^�Q�Хtq����C��w;�.�B�	NӐ}V������2Xޯ��[X	�0f�<����;Y2F�H��/!��@dOs��	;��2�$J9����5:�y]W� ���Ŕ��?���%j
_,}\�1zu��А�u`����+��r�n�ts��p2��Qw*���@Ӊ�A�/�F����Qj[��λX����(U^�G`{�6�
��aȠI٨_��SDU���L/4��HPo�R!�uexj�����H�J��שs�(�Haj�J�H�ׁ���Ђƕ��ڣ]�~U ������ dy����y�
�$�yE[��U��������]p\r����D���6�^�w��a9O�����0n��s�n�W�����dϛ9$`a��'���10\C��A�5,�T�0�H�(X޼�V���nFh��2 ���w��
$t4�1f�M?�M�I���N$��暔�������-D`5���q����ĭf�K	O��So��G.����i�=�y��nR*� �f�l�X�-�E�3�g�Q�rzX1�lfMH�\p�j�����L�PH�3���6XC8��t�N�U�ݗ�[ؾ��G���@S���;<%)��UB�ˌ�S�F�Iv(��\.���NXa�9�K2�����	�aZ�Z����3q�%~�' �l��=8u�Ϻ&M���#��8��#ɴ�w����L�gb��V�T��5QY<=�<:ȍ�Z@�*��B�5�	� (?� � |�".� �^u4Z���'����e�I)�Ni��}�tB:��8�O�5^_�i�����{Tu}�@/�?�}�"�O��9�g�$�Í2J�l�M��:c�W\H"�z_*��N�u���J	�Tz�	顯���؜�ځ�}��Q��R�~�i-flk6D_�����O{��[7	Ј�X�t����<����5fP]����B�u����m���"��Rl�'Ad��vb��c���0��	r����K�ڑ��������]CP�o���1����D���)��~�~��+�?�I0x-֚���:�KV�}��z]:�=Dř�{�[b�齦%����Ӓ���kz��jI�S@1]��(�%UO�U=Q��d��SP7%]���Cq�9Q���c�`E�7l0��/i?Z������ks���pr�Ă=�C{^�CW͘2�٫dQ�(���Wk2��po�)~va��?z���)����>�_$�s��5���ղЀ�g`�`�=H4200J.|F�g��hg��v���ߞo��GK*���� �n�&s�HQ̄�Ti@+s���g�{.���WQ7( ���*�u0B��!����w�����}6�m�I�;����^��ػ���^[{CW9�a��'�{�砹���ġ7��K\L�+�j�����]͍l�i�	̧!�<$Mm����t֜����n!�t�ܢߎFQ��6x���4$�����z��Y)�k�-G�D����hS��2s˷P�;��p�0�%ɪv��2�j}���:D�������jO&�ޟ�M6����{>`u-C �Lh���W�Xh�_6��x����L����*�K)�'ZcNo����KLP�z�6ð����}G`<ecu����/Az�Q
�������
��B�I���_��Pڢ��l ^P|�zґ��֧!�v�l���f���N�vk"��Χ�c迥�42�3��%R���H'�4&`��w�[�Z��&^_3ȱ��i	�}~��m�M~4��H�M�(t������+R{�WHb4�:.u Ju��?�5�ې�ϡ�ms�zy��m�Q�"j� qd�i4��L��_f!A<[�)R@ŋSa�$���}�6�h:C�l���H��Qt����lwf���g4�̽g�h���rZ��v	���+U0=�H9�@Qw꼩e��` d��L�ËH��o#H&������D�:d����t{ߪ��N"��1�5"�½�:d�V��Zҵ�M�%��V؛_˳?�i�+�¬͕〭d���Y_1��#`lW�W����`NGj���揻`rkW���5*��I5���Ї���xT#�5E�׺�sɢ�[;E�N����3�U�~ю�v$���2�Ȟ�d�yP��5b÷��I�hٮ����4?��&�%cm�
?��0����z�3
�?�;�ղ2�b* xh���!��?�sRJn;��7*��oz�@`@팺��{�Y��x~
I<�L���l)&^f�hǛ�E���+6�0&�s��V������Ϸ���x���=^fd�/ -�Je�]J,콨z՞�&z�7I����]���$`��pb�I�*^(�m�^�cRz*��a4�f�����	��Ţ���������7+�~^��DK�'��:P����,�{��!0~�N*�j�c[�*�ִ�qj�#�%�anj�Io8xT/n��0 C/�4@��}�o����V�!&T
�˸�Wڋ����¤�`�䧸2���V���ξ��8���G���s���2,���v�����c1,on�RDe�U̜Ro/�QZ�J�sU?*J���&�K�Z�)�H����Ԯ~/sT� �`����'��L��E�\K������[J��{�}���yP�n�qL�ހ�)���6��:����wB��S�� �RX^�M����i�Nji�D��G��I�t4ܧgc泟T��H�;��KZ�A��oK��_���Sh��:�\�j�ӽ���F���u��T��}�8��!(%Dw��� ��MV\we��P#4Å����X U'�)�E�y(լTQ�������J���ĸE}R� �;R����}b����Mf�7SJhezoB�nk���"�!Svq@�����~�C�������HRj�R�WÝ<��qn��ѵQ
������]M�?S�Ȝ8�����v�gA�s�����1�Da��0�M��٦��֠L,�'*����,�')��8�I�7�A�ϼ�� �8�XEVϟ�nJ���D��l��"�zg�ᄽ�4!�!��n�IV݉n����$+`��V�1m�[�ʸ�wG����*�Yg#K�i�!����yeU:ga<��:!P+Z�˙�4� ƅ�