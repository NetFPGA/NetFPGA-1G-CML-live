XlxV64EB    168b     8b0lV+Ceɬ��rx�eIq8�_:Ad���ka&�j!��m�RY�0#+���B3���M&�2qh�k��t�'��N0v�^#�C��(��`�;7�'�-��@"mf�23��Xuc����]�i�#G�rm����$�ݯ���W��0�ZKP��c��^�}8&V��c .�`{��US�����Q�(sf�'�%J�}w���;!���ul�ZW�f����|JG�y��T�Ѕ���%��v�4��B���_��:��2����Dz��u����0.���W(TQ��߆+���eT�o��/��{_�@Ҝ�_�y-u�,
�1'��E:�Px��p�v48����=#~�=��SHc)�ƛ�&w � ��&��|r3J�-�1�d� ����g��Ņ.-Ą��H�5��H1,f3���ՑPl��\�Y��l�i��3DF���4��.�A�!n��gf0��\\aш.�,t&�<.��)X<�6;}߭�T`g%��ٽz%�y=yt��(�kim�0Q�]��,��>S�`tH��3�Ha�8�t�z@�ŗ	�,-D��l�h����UI|fGZB$��G��>9_��*^N n��Mp���˗����,1�,[2�3[r�[�&D����<������m���:�g	<-MȾe���X�I�\� S%I�%����6]�|Rkް�S�P�lĐ����QC�IpC�M�N�{��l�u��:W.���f��������L�-5�z�"�]^���(��1r���iԈ6F1���Ϧ��MB����! t�~�V�N��k=R�0V�L/� �=r�5���az��4!�e/�kl~>=͈_(1#��ɭ�+otb)W�@?�U5I�ޣ���
�m93�9�l�N<:δO��n��0�X-�U^#k��hi�=W��h���!��E�FA�BH�`�_L�r�hb�~��Ǌ�gZ���}y�K�(��<��Z�+O������@~y�͑"���ઌ;�S�.Tx�C�e�3q����S�3rB;�����P�����!�s����V����і%�t���*����s��B8l���'U5z�U	�aa�}l�J^	 �������T��8A����%o�ݿ\�( G�s���m�F�u�Ʒ@����7r� C�(��N�ԇ�^Hpl
��0	C����P��@4L�l��0��􌓙s�\)���ۮ5��=u�/=�dLހ��+�����X?H�#�;��FI���[*@0t�TU�.�4�y:#|��U������vݡ���4������0�1����"�qq��[m���*�(נ?q��r׍K8ٴXQޜ�e�r�G���]e�d@�D�O�3f�e��b\D;�(�Cϒb����LM�FM��Q_��Q�e���t�a{T%��J���&��~���5�2{���Ʀ�G9�(��5��ߜ流��2��_4��dx����|� T$O?����54vc/tJ1k�A�_n��(eS��SZ���M�7X#���_;V[>��^�+.�y?9?Z7?'i�*c�S�T��"�kяH�Xġ$�`"Uٝ=��wT|p��t��4T��q	�^�K�.��b����#=���LϿO~�k�?)9u�Z񥉪
R�Ѡb��PX���30���ӁF�I)�V�-a�����2�7�̾^�OE��$��Cw议X��j'�=�v�l=LTd�8��Qu���U3�F�c}�� �SިM�sVY�_��[�c6w���6��n�TO�m�P~������4��������f�h����	��6��\,�s�6˔N���Ƕ{b9~]y�$����i¹Et>_�~Uw�ӿoK�w��_6�8�Z���2T2v@�kZ�)�x�춪��j;�q+�8�p�P�X;_�{�L�j����*/j_F#A� ������g�$Si��r�!%E0�}Zi�.5�/�:c��Ӝ����(Y�<z�~�l��G=�l*>��z����zۄ���u��V��0���c�.����J����27l+��]mP�Jm��\��}�jAR�n^�D��3��y�f��>�a�<t�*���(-y�����;G˒o9�6��B#%=��Q`�B�P�%_f�\�k�fOF��+��kDi�P��Y�/���l�4ɋ�%(!��B�,�,����^���PxTmF��͊���7����)�@�H��S��������Y�x)�x�g����