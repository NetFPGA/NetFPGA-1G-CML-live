XlxV64EB    2837     cd0�P�� �W���At�@Ņ�7��q����'E-��G���2�B��fR�����c-e��n�������h@_��~�W�n��{��ƯǗ�򏀷i_�`�d��^܍�	�r�(��%8�H���/��0o̺�i�Qq}��a��֒E��L�	U����TE����N�xA�oZ)�Ug�gNQ�^p�`qk�Zp鬤�ݍe�FdW���Ȁ�h1w8���}$��5a���[�"V����S��J�y���MdFLnl�.e����_X\�
�.��1z���B�tJa^�7J;���Ϻ��p�2��a! ���.�.�h�U&o ��M�2|v�5���:�ٿ�_3h�+@�"fD�~��ԍ���)�Ӿq�M�N�8������T�9�U��jS!m[�;5��G�*��Wd��-�@"�fSo��h���&-�RU��,�����_�meM�XH�r�Ә��-t�
�/x� F�yՌP�Ƽ�8�9k+75b?	�Fi��-���m�ܦX�[��V��ND�����c~���	@�׮��
�[ň??�P�WR4�s�6�(�:u�����\��U|�I^��e�����f*ʼ��[����J��8��7�0nb=HZL��F#���)D!0�OPc��mQ^��9ޗ��g�ެ\��}�}{M^�F���\K�z�)��k�J�H_^����ۤ��
��d�'
_5���c�W��d�JNg��+wNT[D�j��'��1��ț�,�8�̑��-��uQ+���&C;��(̓�<в�^З/�?�ڼ�	Z�� �+�ٞۗS��f�v�i���8 �g�釹�{��pEt�L��#��.����JQ4"�>�O*ru5WVC&�u|t�wD���Bz�����M�@+���tZ4��1X@>��%l�îϓ, �Л�G�=��\R�͍M×ǔ5�t�#���c��5H���YgN�H��1w9��[���}E	�@i8��
qQB7��)��YUk.�o��iUT�89�a��Hn�R/eh�iW�m��u���t0`?�c{����ޤ��\#l��f5��?���?�RH��%�;q�BU�Ȩ����K�SM��'�o.��lsD)�W�乣��~tlաeMLl�4g2�O�j�Y<F�])rM�D���8�f�4�8;� X3H�n|ٗ�/=��)�?����K������"`�κ-#�]����ń�|����C�� �W�wNӂ��P�鴴�;��=��" �Gn5�ն5i�	��>��C̮����p��+q�$��*�
�3�[�Wa�h�@�h������Mg�d������k80`rW|C�L*@d��P���a���Z�)�DE�JMމ�ބ����x�q������d�v�E�3UW^����|vP�*Bݯ���)�Zf�\�D�ұ#T0a�'L���Q�N����_"�ܓ�L�ag�����	p��`=�_�:��~��	�q�H�P-�+�׽��'O��$M��n�/%%�n��>�u t�=��hQ�9�[�yO��y�ʍ�G�ى�暦�H"��yh;��5�?HO���z���4տ�9���%�_1�V������FL"� �WRL����&D!�<}ƌ�aC<r��ME�P�.��s3V�2�T�*����IQ��x�[��3�Uq�4_B;�fEI��j0_(A�͠��W���)�vB��&�T����=fZ�ͼ�������Ք��l%I�^T��GK�SoC�ƭ��&�dx?B�~���������]��^�G�4,�[��ߑ�5`�ݤ�r��y]f���v}c! ���"km��e���R`��Z��S4�c���fT߉�?���+l�
�����ɤ�q%И\�ѭxe����jy2e���ַ�j�)&�-P9���v���&`_�U��GIs�.�
-�ϰ�PM��H
�o~��Rׂ;��z4��O7����Q�]�%�z=��e?�UBna����] .��..����->��;{_:a�y=0��[�0�������W����$�G�.���OQ��6�J�]C�蓬�s+��H.d�b�
���R9-�w��n�tI�RZǇ�#У�˨��g*����Cn�qV��
ډEѻ�P��l��*��躾��z�-D����(���fW��<�+���Z�\�1R���G�;A����Bs�	{�	�kYy@��}�!��U�v�����q{� ��,<����Ƨ%o���F��%�St?�����k�QV+z�'D����.�=�n �������$9+2{���}~gy�?N"a�h�P�I�a/�����m�
�!�B�r����Ɗ��Kϟ�DvxO��Z�y+ͦY
f������`%Ed��w��sţ��Ab��X���@�l3�SH�לB��ח�F�4[6$lOƯE���˖&�V5u�����"u �J� �Hԡ!��B�7)��,E����-%a��A��¹�9f��8IjĹ!2��Q;P�M��$�z������wޘ:2~p+8���)�Q`�����8��2�]���`Tc�����d��l������7(D�A%9��O�mӈ�O�!sY�D=>1�|������	$��ʚ"��n�8�^qz��Y�$׆�lNB�lv�m�d�3�F �a:�[
�'g�b�uS���B��J9��"�@�zg��_�(��Fy��R K����j���򑘍_���5�gYQdڐ�c�-�[=��L�I	��e��.m��&��X��f�DT�Q�/�ݞ)T,[^�(�D1�+�6䯨�:ΰ8����["�jv�;��K�~w�=o�qF��c�-z����g �Z��2;�L��i���?W�R�.�W���'E̗�K8��Ր�b��R|����6�"Ƃ�r��5*�ȅe��J��7�%����0����/=� ~+Ɉ�R��.։27��8Ae�xNj&�S�|C(c��t�f�x_A_�Ӓ�U7�P��c��Jw+��ѹ�����H
�-D�E��������R�v�hҭ�	���xp^��9��Z@���&�q�W�kc��&;e��O��Y�jT�f���'pq3�TɨQO�C-��~�˦:cӕ����JX{���"�e���[�wd1U�rJV���^�M|w����Q���x<gK A+�����@�v��)Bx
i��SϨ����y}UCFi=���V�;i���X�hf�
�