XlxV64EB    1feb     ae03C5�?�����2��C&���L�텇��|Z�0h�%搮"�pE��n7SqȆ�h���&1�*�7b�?Ǩ�,����G(oh���q�g�v��T��ЦGJ$2��k��w������"���r�:���nD�
��a���_Y�������b�K���� V���{�N4����e �܃�8���$��U�G+��l?q���2�ކ���Gi�����ś�&4c����8,��<��m����fg!�&dX�tbI��X���EE�2�v�f܆��:�iؠ	(�{��wh���*�l3m�L�3a�V��J@>��X�Wɒx49�I��@-0��&AEY�H��ƌ��޹δ),}����<ou�f��5��#�i!�8��6 ;����o��'CAM�9�ǃywN���n��f��{��CUӮí�P'�l��PE�+sP, �����-�X��c��w^U�m��ҘKxB����?�8k�:��u�}x��o��~���}!0��e�+��B�?y*�	[q�K�e]Z����Sk !cL��'���7�Xc�%v�~��IX��_�{3B��H�F,�ڞ{��y���m��OKs������f��;��}�I�����b\Kc���d��K#�	#q�վ]aSx�{7�N�j}�D�g~�_>��:��!Ȏ��WV\�j���z�47��.Z�ދ<���2Uݨ⩕Yah�7����!�I��S�R��Iv�h��7�]W4��W������Z�D��څ�s~yB0�t�}��T��.-�牱�_`�K�χ�$��*�9��7p0M�4����1wO����=��T����tc���v�����c��,����{��7W8O�,+�t�?�-7#��=IX�D�����^��
"�ιL�!��晛.���{��2�B.�d˥]?ޖ�4[����b	�y$"P������a��e�F!ac�L m�:\F<�ߌ\a����	KJ��S���zYsb�++�3���|��罽y�ܦ�q�L���� ��qL/�E�VM
�(2H6�ν`��H!t'~�k��NI� �s�?��Zt
]�J��������'ɕ0~��"�Q����t��Y�.���b���>�}^��Y���?l�Hr}N�о��1��-&6dII����P�ˏw��W?�����3r�6Zkc�I�W;-v4���8���o��YoU{=��>����@�y�K�m�����t�G�`�g�8-+�\P��u��"�[�[�W8����Z��=��b��Y3=�����m���yn l> F�k�rN�#�R��C�E�-W~�z��Y��!a�j)�/h�jL>O���tE.�J���E֯f�)�g�T�޴��t�����Mcj�)��Wuص��V�dO��W����pHc{A�XN舲['�?lfi:5��b����O��_��ŗ���r��|b7�w��v�%v}��a-Qk<W�-��9X�v����p� c�3��}�%�Q��7x{]��<ҝ�W��q��i�mP�
D9�?Zƾ�i/e��1�d��25@��f��՟1ْ�D�7�뜽�����wz��ѥ���n�F�ԀM�+:ְ����W/4h�Z��z[K�f�,�i'�L�)�"a�۸�_2�f�}�c�Y�+{G�<l���P�U�P�n�������t���	OΛ��� �u�
k��������,#��>����C��t�>�y�ѐ-y�P5�G�������_:�ʯ-��Ik65̓}�\G'O$�T?T��S�[�̘�x}{�����Ę�4홹�H\��Fy�b��]
ߢ�w#���'L��oå?v~ё����$?1k���M�]$�b޾��z_�1-�@�2Gc.JM<t���������������s�_��8T�H�V��<�(�(����H��V���t�ž踚f�2�y�}U���5To��3�{k�As�m�,��e=�O�=�����
���n);2��A:X��l��2��(�l��9�G����ءL���WT=�R'�Z�q�#����X�	h6�/b����U�1J�c�����4�MDm���l�kϢ���H&�BHe?؝��x��#�?���ݡo��?>�孪�8�r���%��)Rj�@��������uk�A�k��I&9z��/c����Y��?.�R�O:O�}�w�ut�!4��"��@�K�C�Um�q��40z��ͣծ���b���Ɔ�hČ�v�m���^���ՉtQ���{O<q��_��}����W�ъ�:L�϶�'�[���Z�|B�e��b^>�|�`��,�:uz���'mr�%؏mA�2ON��V�C��?���f���m�
�#��Τ�8����3�氻�.)���~3���bY��}[-<���yn�%�j��C��KM��/�DS?_�\@�6���1<g�)Lą)2d�$L=d)4%=��⃑���i�����Bj�6Wd8��_�ri4�;�<�(���߄B��D�IB�
�'�<��D+S�o�E�L$B���ra����㯮����Q�����i�l�m̑Y:/�+5��o3с�vM��8��"E�є�v�*:(miY�if���ݳ����0�+�S��(�ktY���4"2�>�z,�/��c�ȉV�N�k ��oM�n���;9���Z�`��0:N��4�oԬ�~�b�� �� �;�:�6-\���[h�