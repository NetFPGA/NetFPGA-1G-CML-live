XlxV64EB    1573     870�a�oQ5��x�k�%]���U!oPx25��͒�<�[vb��q��b�a��b1dZ��J��d��*�q��K���U��b6�a2�@��79���@�0+��Kd�7�D kdf�[.x��è����\���/T��	����ԥ>���rPpV<���n>ˆȂ7Nײ�B͖�q���2�gB+�C��G��,�y��{�7@ڥ�t��[���u}8X�r��!�a�yj'X~�v�=O�A]M�M�Tvf�Ͷu$��������t��2
���D�W��Ru�Z���?Mu5�(b0�"֜��.��S�d�)����v�߮��g*����}�
�D�$\:���)ȃ��+u�����2���QP5~���h��qc�Q"h2���(���N������L���u�`��T�nز��̠
�8ON�i��E���5Yu[F��茶�E�C�(�3��;9(F�ȭ-Se>J���6�����Q�Vo�7��EP+){}�c�m ��^�g"��Z&����+4�W!=�oZR?�D�O+�cg�5a1�����hQ�y��E0�m���B,�_x�陂�8Bc脥��a�Hav\�t䅉 �)�B@/,���T!�8��"�³K]�M�_��V�&�	�/��Y�8܊��#����1c
�D�:�\����W�Qv���αH-��}y(�Ѓ��$��F�+X�1+�-���t���׻e���]���i��;	"`��f�1b��7��prs�Ȱq}qN�!�N?7\��e�t��l����_��b��c��,�	�49=����F7�p�ԑ Kv��a�/^_��}�M��pը�߶&��d�H��������G�9!z�Jڕ*��E~��|�����k�)�=�i�¬��_�f�E^���4�a�|v䐕������>���~_r�_V$R�&
@�1F��t�0l7gY9��;N����P�����c��c޳j�$r/n���08��X@�OQ*e$nlו��h����Ŧh���8.�F�u#�K.ANg�Ͳ`�9J�Xt�I��/��Ԡ<�"��QE�F��/�rL�"d�cc��������Y�4צ����u���"�Y�a0f�oC�j����k���'}D?P����c7�f�/GS��s&�O�1Yc�奮eג�W]��i��Ķu"��p'������Yn�&�O!%%:|g.3��O����KCu��p`ϒF��@Ez`����eR��5�i�F���ԩNWy����Z	���R�CA����2�)?z�����ĥuw{�a�%�MN��+`/��@b��f�:td�Z^�e�}<���+�O}2{�SDzub�dizm��5}�D*���{��q7��᥁��L�Ǝ���A��~�Y ���=)3g۪���
W��R+dr��l$�����K���4��9!8 ��$a��nC,Q�ׯ`��:���s����Ϝ�I����w15�񅧸"Ȫd̻�7\g��yS7A�H0ܸ�;�j	�[�Mi�Uf�f��{ 27�MJ�9��y
���$;Bn�f������!�N_�;���_�I����
�Ht�b��
�H}��tx��z��/) ��Q��ӻ�Jۋ���^T�&GI����t��n@>:�<օFL�
�5�����i N7@U|8ƃ(��h�:�6e��� 6��-3Тi��#`�c�P���׀�Bح���hT�����	�]�xa&��i9�՘�woq�!=����ú�RY"��5:8��P�N۲RS�܁kR�vuC����y�(�U�HL�ު5�?bc��Rt��9n�S�2�f]n'n�qS u��	8(��� ]k�@�K;����Y��;�%�U���@��XEJ:~�+C���b��h�[Z3>p�a�M}�%��P�jES��$��yo"k9��T!����0u����-%�U�4�#�5µq�[���)��RhuP����ۅ�oIY�A3Rʪ�?G]h�)��3����6������f���!(���I���n�4�;fi�E���aܹ�x��^����G���P����B�Z�tnr'\�s'{�B��:m$�ke��Br�*J�,J�ʻ��l�߽Į����9� *�؏ޝ���=��u�+�,���