XlxV64EB    3203     de0�I�u�S Yw9���UFI�C�Y���I*pl7g�M;=g�5cE(�ب��o�W�?���f!אG8���Q�o:���%��B'
�G�ݔ8^���u �`��|��YOv<�7k�o(�.���횐"nhe�0&�e�6�,_)��^�qN'��a�뎴��ف�7�s�Jc���U�c���z�ך�r.ܮ����AK�}�	�$qߚ~E��b&��?�S���s<�D�jU#�Y Љ�d/�[lK[ߓQ������ie��k����{�o-�[+���>��c�8��tz\��w�Q���hI�&2�`��q�O[Bo���,D��gL�jfzir�	���]V(�?�����% ��?LǷ�Sr(�o��m� 0�#q/����(��lq}l΋�2˅�nJ�ޗN�}b���f�1�fF��?�$.�!���%���/)��2���T~(���g�;�"&���T1�k^Ζ��%r��/C}b#Ox��x-�/5t�_�v1�]r�-����΂ �ۯ$�	�M��5�3�T�DbZ�"�G3l��tg�/h��٫�]�>Z�hy�,��[v�z��	���7	��.�A��H�_B����B`D�si�Yζ�7�is���}2^=#E�� @�G�����í�av+��2#[�?���� ��j=���Y�&�6'�T��ݰ��!��G&_� ��r���e����L̦��R��d�����9�k�%-�Rf�R�Jj09H�?�b,�J�8���9&H�����ׄX� �8��Y��9��7� ����սR�Xj� :���/sy��W�ч;g6t�6�?R���|���=Q��i���T!��:2��Ҥυm�	�]B��D��i��N5�:]��#_���$
����Y��
j�	<������*�+Q��_��^����0�O���Ε�1�����
:�m���C�!��}%Ɂ9pH�!-$0��w�y ��k�>�~��W�w�����4�<���;Q��{m���d>�H3o����Ѹ�0�\�J(:��B��=�)�$��+�E�k�g�jdG���ys����mK�k���e�ٔnfK+��d���ۦ������OZб]�'ltG���*�}�d�/
g�@ں�x#��çE���'Z6͙���[=��R���z�������� �`���7oT�����Xʚ9;�`�4H��he�v��3���[T&��	s�iĒ���g���2�;Z՛-�>E��:M���Wk��qj��h��d�d�б�l�~R��{Is�����]4@m���q��^9�������:��綏��pg�8">���!���Ϗč��hz�W4�sAhnX���R�m0�º?{#��9�Sz���]/"�Z�J�	��Я���#iM��~�'OYl7�B��
LCS�B	�b�S��KId��v�������K d�c���?�_�������L�_'G
�cy�����}y��q�#:�T�X��ĊxB��AG�����t�F,%�b��m��_�w������-,JFNg�<�}6_�I��l�go�rez΄s)�G�)�����K��}��h�$�F҄�?���!�-�Q$����wM�p7Kt���� Yk�;d[j�����}H��ߘ)�h�jp*�����]Yn�O 3�ǑB�h���%�p��|q�.�x&�c+�zn@�S�u�x=+����컋��ShZ,��@��4�����(��/��N�sK#�?��$��΁wO�q	��&���`��9�vZ�m��Bk`�b��d��[0�wI�.��ɤ�gOl����jaGj��\5��(1;�u�p2O�DV4?�*l��ׂ��t�!���������_KhЅ���qi�m�drw�Y�ɝ��;O���J���
�(�9>j���5/>�~�Թ���*j;����M�,ÿ�oHy�&$��m���O~�3O<?��7�:�-=��}B���BQ�����HmĲ���T�&�y��1X`��6�U ֍T(kթ!�ن_�����>UUH�G�?Cy�O�"a���R�S�l��k�b0b���^�֦Bī�1�*�d��h�0p�h&��	�j�z�r�+l��̥8�w�)�(~� HÚnV&ۨ��~ܰ�ķJ��m�C��o��-Y�u��ٷ2'|ê����:��C:����"	U����r_٠h7�Uw�*����13A��o6F["�ޭ��[�G��Ǜ��O9��K�0���@7���:����!S@�4`:�����>Η�����[�c�u�8M��؟��S�G+�9KohE�q	C���3���|�H�]��9j�������-a+��-�VW'��^����r/���	o��7�I���4Q�7���ޔ<�pcz
'.)�7�K��g�Wm�!B��*��z�"ڢ�@X�E������#������	gw�}�ck:���L�K?����+=�!��yqy�m���쇺D8"��f�w���wrq�E��h��`��%K
&�dчޞߎ���V�����h�+T�g�U���G2Ad%�� 8�|���jA�f�)�������b�^��L�md\R�.n�%��`�v�)"&zp��|4Q-�މO
[O�)�Uh<A�`��(16A�1�-�A)�:J�EIn�=h^��%�����T�ϯɷ8�,!Ck"*y�%�ļs��~��>���'/1��-�ɣTT��DbV���G/�z!O	��W�Q"P�EL5ij� x�Q<
?k	J�g՗XzC��n��D���a��q�~g���#�S�^��DI��U���)��s���l����mjC/�e/.-�Y4Zb��j{��#�w�Lo
�4Ҧk$m��_=��]*���Nv�׿X)�\a�Q��.Yigll�>s_���xn'J����I���6�!ۘ��bCl_cU��<a*4�jR��D�k���j������C�ux��W,��<-�qt�V��k��FQY���-�G/X@"�[9�}̜���G���g^�1�CU �!��Ӧ�R.C��\��������Ï��L����KD=⩽m(C��Y&�A��\q��}���j����+�
3���OO��'��8��V��*�Z����0����a��"�;5t�iW��i�*���B+1XSfSP����u�p�ك�z�%+R2�}���Է��OG���zM�Z������$QGD��4v8�X���ү���a�!E���齶|����]H��sp�i@\o��N���|�*N�hw�2U��|����ju ���p����X%�|����	��k�Vf���O�Y�:��(2�W��n�i3.���`U��|��`�[���Kt�x����Z�QT�.h%h��5'MI��u��%�����)���;�2�H����Ui� +�#�N/�ӳ�r���ϙR(`��F�.�(W�g1޽����k{2�Ϙ�jQ���^�ur�&�Le��XS�f�׈��[I刖?��d�<ҩd|�>�[�����0