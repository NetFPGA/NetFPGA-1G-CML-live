XlxV64EB    a725    1bd0�v>Y��.j`?�ͩ�������NP���K7�+^��3��*�f��f��r�K�o7Ř��X ����p��ŋmW ��H���s>W��M�He��<��바���`ё�� r;�����ao5��E,"�k����[���,��Ì�o]��`A�k���1Ҧ	��m�GgO���9�x2�8�ܐ�u��D�.M�ļ`vs��4p�\����b����y��z�&�b* %.Bsg!S�lk�T��Z\�9i7��rqݡ�@��2*/f�#O�9��l��:��ޣ�]�?$me�nݓI���i$1�L�!����^DlM�`�jh�l����ɧr�Z�!�1HI�բ�mM:ڿ�H�4���9\4�W�
t�Uz,D0wkA����̈́+L[f<e��t���'�8]4[�00f�r���2�p#�lM��=&5�^�O��G?t������<;�t�:���2� ��rdS��z��>�Z��Y�@��]�'�������n%`���<��.��q��L��VhQ�~�J)j�B����3b&9�U�hW/)�i�әV7�ɘ�aƎ(�da�$ `0��s�1[	�<.WQ|�CHq�	�q?��(î�I7W��� �{
[s�F£�@�#v0�Xs��6��Qu�yz�2V�!{�OS�gN�dQ���s���\53P�����~S����ʨXz��^��]�9[�Mt:?�}����HB�t[���-�H��L�Zq���H����꧰�62�'ܽ���idW�'���*%�[��|i��QV�<5Ћt���?+�Q�G��[LTv�2h�:E*�ڪ	�� Jp���s�̙����?��fe�cb_�3&2yk�������/;����u�9N�$���լj�8�V ����~S��O1�~$�b�?�i��P�>��0>��?qڧ@�����}�$����)�i��Һ�$��Y5Ϥŷ݌���b�F^ϒX�	���LzK�v��=q�ib��v������;xM��;����=�vQ/��n̹g6g��f
Fzu�ݺ�X��}�wU�����צ�3)����'96�*� {Hx][-bvj�V��2m�*:p��<P�?�r����	aŗ�B��V"�J���%�d�:�h�&�t�pǕPkua������߳���H���^8��\���g#�+V�D�z6��(��/V~���&VO���~q��s������1����������zO��g�5������L��O�9b֒2ڋ��N��^�h*Y���_�e
	k+��c$��	�N%ۇ=&C��S�V"�D��<�t�A����\�n�~)��V�{�k+��H�c�d�:axv;��E��8D8!҆�/��[�y����v�W��o&6�5�}�4�
�Ҹ{��V���I���YŶ̊T�9l!9~8�Πb�Y�M�r�v�s���AA�%�awJ�8���I���6xP���!�_��u��&�G&8fW�2\f���?���\Ww�ªa�36��� ��:Ray�H�u�a��О}���5����1�証f ~�/C&�%0e{=z�&a���C�2b8g��ޏ�� �L���6L�V`����'Uǉ�W{�o����
h,.������A�\}�
�eˉ� ������[��6�Y�3�7�hAsJ�6�l�C1T_2w����駎������q&O ��y���8j-����t�[��荄C�T�Y�A���o|� �@��I!k�3ć��m?1�IZS�xp׃�Pp?��^�hP���pTBB�e\�P0&t���=(=؁� �]�w||�/l���#b"?�U]E,�3�.��2X#�6�K�[�)M�V|�����:ۏ����<y�Y��k�a�	�� ��Հ3�=e�J�'�������8��z�K�^�W8
D��#�X1��ͮ8�9t�_!��)�*��Y7+y;���a����W�[rE�Dz�|��&�$_�b�e��$�ZR�d�`�[X�vSI��g�^�Q���Z��0k�.��Vk���':+�˫[��I�9�v��K��f�e�ySdն2��~P>��g�<V�S�p?^2l��]rDW���	7�\��IM� �4���~��޽8g�bi\<��_zr2dʈ6�\��R�~.椋+�0�),���P��g�r��5l�g,��c�:�M	����ȋp'��w�JuA����˜���=$l4d~���Ǉ�^���*ce�1Q������%R�����i��ܕ�	U���ulZ\7$�m��أ`��c������(ND�����f�U�l�/(6JJ�R�ۖiנ@Ѥ/'Ԓ��#���)EͿƢ4$&�B��T蕦�P�7����)�2S2w��rE�GA v����&� �����X���� wEǕ���7qA��`�g�����%^�#g1)����`�}��O'8:�c�o��M3�����[��(A����ɨ��ڀ��w�G%#�^�A��l�r3ؖXu�'Dj�� ��a�%����xNNǡ-�¹�ʹ�,��p.}Tj�^�`���vM{T�9VFC5�Y��s��/w�����X�
�WF��n�A�9^��k\���&E�?��Y:�t��ߌ4�i����~jO���c��l�u���f��4;�n\k�R&-K&0�:T=u��/�B�WTn�晪��]��B0OՅ�o�P�����7и2������� ��/Ⳟ�2��[d?A3��.����F<5�5���j�D}�O�/UP5~��jߣ�=@��k>�H[[_�.�]��*�L�g�/ �m�z�ݱ���:ĖlS�I8{r�>��8���BcY��ꒁX-n���j2�ל���L�~��[�M��]��gC���gOK&��,�=n����9h�[��(>���O��F�o���3}�)�%	�kc`?rIx�'�d
&��]����M����̡u&YPS�����m�k��c;;b��;�я0��
)1�V��^Lx��w�/M��A�x>X��nDq(�B�u������ue�x%-
�����:v�9Ӛ�C�J閏��y���*��2����e��|�6L� �ź�|��\+�	o���9y臗�� w��ߗ{�g:��I�T��
�F��0E�����W�i�ɢ�\�e���B��aAi�nc�N���+��ǅO�E>���T��0<� �3�sV�Y!���5�(�ƻȦ�b��ʞ�Y�h��k�7�4q�}	f�ȸz�-�6+������,�8S���t:�z:F�V���?Z!wV�}�S�G�!�-"���P7��rD��&-�H��D7��<�3{��aѺB,��o��g�ҹS�B��+*%M�m�,�"� 6jN�i��f���>��͗d�e|�Z�����S˴�F����;T��d[�l���g��8f[����-4�� 3kxډ0�D�R-�py�O}�R?_��V������C{ȼ���o�6�Z6�y�i*���`En�LMf��!pܪ�������	/�0������y~i�!�|��n�nI��; 2 ��G�үQy��[f��S�:L1�.g�wS���&�j=�W��pN	�������G����i�)�2UV� ;��ު���-b=��F�s�G2�)�<ho#� ���Dv���g���۴S@[�L�	�w���ń�i 3T$m���S��\����>Q�z�R{�G���{ݾ3|�*�x)��?C}c��}n�_��$ŋ��=��,#�=lޏ�<�ܨ��e������7��8�b�;5�j����-|�"�DLe�;\���Ǳ���io�r���{5�����ײ#R��Ų�έE��� ����m���+�F|��"k0�9,�콖^Xl�W�Ɠ��I�S�Y��M�G����U��}vo���YvKz��Kϟ�s*4����h�
��&��������92���/zB���<gXTeh�*�&Mv�OY��h |76\%�`S'c�&�D/QO��K�j�Yo�?�)�bv�_A��jƸ��:cR�f��v��=l	��,�0��A����CJ�}�T+/����+�0����@��_��x�G5�xzcĠ��c����j��D�����ͽj��,��%�g%�;uPX=�A`���Ɏ<g��C�XI<E+���؅��qȷ��������K�Dl��4W���>�x'F���u奱fb~^�r|�c� �	g�&*V�E4���Gb>MnRu�0��p�m���JN�o�������dz���c��6ݧ9���L;|�%�5t����y�z�P��U��'Q������a�ۡPݒ�.�6�s�*��uh|���jzI��ޢk�n�7,{p)t���۶��B��}139R�
�^��~;W���*n���Q3����i��H���R��l�O�z�B��2Z�� �s^��J��U���}e,?6�-}�	�^�Y�?(&���K;rm��Q�*N�E�a�qB��2�������V�����z7|'<-F�y#�7�%FM}�&�Ȭ)$�2�����w?3��NhM�`���c<�����oGU��ߠy�Hi��W1{�C�n��}��٬��Fu�eID�.��-��Z\��Klӄ�3��B%�4�< �t-_��I?��t\�%:�C��l9{���է	^?vq��$l�}��w�x�JF�����1��xG��tG�/j��x:���A�T�3ucw����W���9/��NFu�Z���z������p����#_JŊ����"&�IV8O��P��Z�(�R�u�&�_,�.��$z���Y��ӂu��O��~�QpE�WK�.���(�������g{�QH\�fj�x���A�|@��y5�Tu��->˒&+C�ᡯ�(�a�Q75	����)�7�����{�~TJb��)?�ś
�=5HF>��k�����B���}���"ye��27K��BRP�\�Оy?��Gr�c�{%ݳAֽ�����Q�=X��A0�thU��i��)�\z�Y�iL8���
�+c�>�q	�hD�dU�/L��V���]�ؘ�K3'a����>2.��] �l�i�V���[�!�p�Z���Ӡ4�𨁩H-��J��'�d>�y�!yW���y)�H�z7|e�@�7�����T�h����W�7-��������]&�%V�ߺS�[ᄀ,px3��-k! �{�K6
��HJ+7{�U	����%��پeR�͟��C~���U�.�����/�mƉwq�J��'�ci��� �=X�)�;ٶw��<���7��mҖ8ps�mL�.L����2 �\3�b�	�&������5�M8[��S�(��eH��GME�C��ᲇL  �$�D!t�a=�q'���/��v!�-`�c��~7��8T������
��H:�{K%�Ҫ]�z�6eE�n�U�.����[
���엀b��7�`��**3��Q;�®�<��J�r�.� p���Ü4�u���rV�(� 
���YZ4��D�BS�%ክ��)�oO}-����,:��}��d�e�?HV�Z��}Ҏ��M�y��G-izM���������k7�ʑ[������}�2�h���[�LF����%��U�B٦�/�~<}�I(�Ul}���y�nh�v}셙���y�1e[�t��|��#�5��=�@�(���l�͝��1w�[��M��S�f� ��9������L��C��x�#g�)׼wνt�d8L>�ݳ���<�ih9�gc�b.;*�,9��|���G_N*���hEP� �J?�Z���j~P]�קM�i�	D<�xz�����dNqf3]4��~���p�B������R�����XHd¹7�fS笰�jh���C�(!.M#4I�=�	�#c�i�8_�y>�M�\|$������G�ԔK�w��Cf�ު���\��Qdh��^��*����d�~ҩ@�D��_�)ݢ�	H��z��&�_N. ��ԓ��ѳ�^��դ��ޣL��m<�� {�c:�d��/��͌���d׀�֨�&���'SC��``6G��c��� ����M� ���>�:ލ�K�.;V�bp���������5�Ƴ�6ޮ05��*zVbp�v@�R[3�h׫�гG�'�����_P��`�������I ����=>]
����9D���V��a�~��Z���&���P��	�7#7@Q�Rǳ�B���EN�|ʨ@��e��$MdD��t�o�BFw1��Z����H�f�`�kY�0��0�j�qmMI9ܒ~���W���!XS�7L*��z���f?��˞�]����S$W���R�_� �A�Ԡ�Og-��YM)�諗y��
����s>s���`I��~�+�|�胉�r�("i���]R�ߌ R>��u$rv����-�#u ����!l50��N��-ݝ� ����~�g5)[��M���_�_��������k��}я<�����z���嬷7׬۵���O�p�K �8�L{��=�(�x�0	O�B�xC3��at�z��&
�P>jAe/U"\+�����`H6�ɬ����A_��I��5+�<Fo�f���Na��s�ɻk�˜jG�]���Y
�ErH��uZ�B��KI_���ւ��}��!ʐ,�2dZb��W��,H0g�`!kr��Yʗv�~����|y)]�j�K�Id�歴���Pu�c 0�WF�C�O�#���A6�	����2.%(����y#H�2�m5��*�<��cl���7�pm/0����QEڵ�PM��#�����qx������y���\���2���3���\h�%�G�Ya'�q������9��7�ρat!F�a� R������1�|����[1������j�X��U�~:2V�}��q���+�;.��|H+���2)���^]����1��WfR�N
�,�lt��P���Ku����&(!pJ�7���ϚwtM�/U@�9�o\�G{%�uȪ����׳ڧ`���W�Ɯe
�p�;D��z