XlxV64EB    1e41     a90RA�H���jF�9�Ih�������N�ωN�����ɌFTp&l@!�̾e"2cTz���s�#6߶�е��@h�RW��-��F0��6oF�hE�XK��	fDDh�ޏ�r~�f!�9��P�����uҺߍ3��J�_F�4h�V���#CŮcY�`O.q���_5 Dj��j_O��u�$Τ�M`;�T�Tx�&$�GH
Fj�%e��D���M���ߤ��]�O��>eޗ���tç�k��iJ}e��L�
��8%��Ltj��b�u���hM�e>�Ac+3d���ܶ~P�1�'f��G�z���m�N��?���ׅN�gNor� �r�T�
�i�o��g8L��X�z8k��Ԙc������لvkyכ���Ʉ�,��+gb��EA���!���6�����޶N���$:����8Q�=��D.�1�g��RE�㍍�{|=&Ok���2J^��Y"���]��.o�`�z�bg��"���rw5@ѿU��(��L��+[�\��U�����_��Q��������ީ�%R��fc�#^p��T�W���&h���kf�1�:�#��Q�.^ioz~Hk��a���[�T�OC��<}��F_�2o_���o��$��kJT�Kg�2x��V#��=��q?sZ_i���hDZҙ2��Q2/���2�k���N��:"=[�dl���Mw��a�PMHmp�T9��d�}���D���X#t����8��]"���}2���)Y��aP@��;-C�S��]?w<�ߋ�ا��T�3�GN �J�bB�o�ZD�.��:
�Dgh����,���@+�[�2���{|~�RW�jqV:�gRI��M��{�h����0%|�0D-|UA�Bwn5�5=}1�rЦ��G�@�q
�p'��b�J���qb鷰p�qj�l�ofA��Q�k(+�n�f$@J�?C�~Ԕ��3���C\9�K��s��dac����@x.������b|F�/�(:���\�م����{��W��P^XI���jI�P �Q9���(�G�:!��{ף`@ �����h�f�	�� u�����s�`�S�3���VL9?�TW�-�1�	��
-�k0E�ڝ�,�,�oe�R�L-=V|��t��M.�T��*D���I��T��`�>�@W�w����I`<T� �;rV�v]�
�2S�	2�@xhb5���}0���a�mf�q�#�8�e}�\nE̘N���>Q��d3d-Vl��?�*�B�����i��	��P�6���$�7�Y�e�W|��{�K��m�+�-�̕&Q�$$c����-���@���o������C�q�s���X�=R�wwG�E`��]�(Z�Ԉ>1�����ZNqa� ��,������W	�9D4�����~o��k�s���5�}f���"��2u)h���֑_EpD��$s�[y����;M�(-�6�
�h.�d�2�«m$�"c�ܝ�U�]�,���z6��b:�gȼ�6�j�(�%6%�����hluZ�ɏ�խb�@q%��]��G0��҉��t��~1�ڜ�{�GA����E����l�#Z��H;�F�K�:�����H�ϕ�KI�9�q3bGܿ˞�a6��͂�Կ��$y>N�S�}��0��f�Ы���$�@Ex���#�Z0Z���%����w>��x��N/�d��]�?k@{��u� B��,g��C��se$���ޢ��ȇ�ԣ�u�����&]P��<�y���O"�`�۝0B]������ތb��&�QL?���4e5wK�W~:s�C	v������tj�Zd���Ev��2��L��nT�́7�vO�DHU��@�F=
6�,��5�'�2��Qi��d�EE��X�њn��w���<�#�i�ݘ����M�/�:	B�鹿�f!"]ԯ�����ޭ,s���������j=���)����,�� �r�&ũEiHChMmXw���/<+G�v�[�����X����m[9�-AY"�Z� �Ֆ���P}~+kr��^�u!iD�#��2r�����^	�Fo�ڏ�Ж�֏����b����dJ���@�ґ�x��� >�X:S�g_S�|P�q���
 -��dU��dA�M+CB�N�B�C�`ՙ�Z���P�˯N.� �P�GF�ٳo�?�t��jB�4�����k?Ń����k/�����Ta(2<c�WKo����^���gj������q������|l�Xt� 3��~+I�������1��ٔ����ͻV���pc���Z�qeg��N���82n��!+��+�hm�{U4�~Ğ2�do}�V���Z#�i���8A��32#sf��߯MPO��(��j�#M��Vk�g	��Y~��ȅD�8�zɀ+���r.���UFPQ	ɻ� Q�%�����r����g�~m�հ�@�Ue�͕�kY�T��m4e	�m�|MBM��Zh�P_&LA^*S=9U�B�`y�n
�2䥩s���#I,*�f"���9����n'�h�K���YN�x5�"�J0W�j���і��1�n(�a '�k����w������5sq|o]������;%Ք$1��þ땷U����#Bj�'Λ	Z�㣿3F��@T��_H@xF�$���J�׽��w�S�K�9%=�p*���6����J