XlxV64EB    6e48    1690�q�\+m��:J�$]$
���ԝ�H�&�����n��}v^��m�v����;l��!�}�߇�m��B���H��7�T�:^3Qu�Wl�̒�B����aר�W׃�$��S�5{؆uæ�:�
���W�;�5���IN���.�\$y�z��bl|�3���W����kC��|2�W��G"���[ﵜ�v7MK��K��Y�v)����nv�o]%�.��?��x��[;�HR��v������}<�SU��k���2Edx��e$�tp������dUS�����6��,��s��
|�0M�Agv1:��w��r��Z�%�Z0
�ջ{�1��0c1��X�5.5HD�M��&$ݣ���_���_Քk>�FO�p6� ��1� ��з�4�-�
(L�T���,Mw�Ƒx������i��_�M
j���Њ��5)���z����@�,K���C��j8�n��J� lQa*4`�.��&ݍ�R��+Gq�z.�J;���	V�~E~��I�O- �q��1�e��m}���ˢ	{ꑣ~K�Ҙ_y��G��`����u��3ױ�}í �@s*�UP��f�笹X��ǡ�x��k��'7�f$��Ţ=�fmG9.?�쓍z�2<�^e�YE��ݤq�ί���Y|J.T��SM�aa����W����ݧ���6��Ė>ŝ��HI=l6�Y	�X9��L��(�b��g���Q���V�#��am�������ǲv���)
��po���Ls��n{rbU�_%{�ne�֚!��`��dD���t/tK&z/H��
��k�1��SB������L�{7���t��(��͗�?�|���݉�c�}s��L����4CH�{2}�<�Q�B��W��@3��J��m_���§�ҳgB_�(�͢,�ac$��_����g �S��l�����k�n!��e�, V23���������.a	�N%���XYd&��aѧ�!���Y��G���^�iQw�Z��屏�7`�9Zǅ�V΀�P���Y��p�7�L���ƈ��`�M+��~�T���������^6Xؽ��QA�d|�!cz*��"7��ee��H�5*�)h,�x�%-�o�`��|�G9��}R"m�c���'M.�{�"D7_��l��'%h[^2�<{L������*ȫi�6Jf�u����[}G��褖�ຠ�~=%���a�8<R�>v��H7� * ��_�;��J�థ�9�S�����|�y�g��4�ï�
C뿞?νm�~�,��	���
��:%sJ����;�m��đ�	٫֫��Ϩ����²:c�QY����2��4 J"w��!�PZk������T=�e�Ζ���{�GʉC��>΢3&%�2��o^����m�1-�%����Iy�k�����#�M
+v�q�j7��Y90��d �+#�/���������{���&���['�v��:#�[Ƹ�t�k2�#�F;�!hxQ$bt`'n�J+�Tf��):*zo�R��f�LBT�Y����,��"�q��A�?avj^(�IU;�I
#��-�Q��%� �z,�uJ�*0�;GȊL�����w�*�,X>N�#���}�=���o��sE��/a</����	�����_�7h������)w�^`k�<ۃb�M�yy�4�'5lJ�I�F <�?��I�������
疌#��� x�DI�ORa�/�Y�Ҏ�m��n�.*��g�Z|6�"�ȭ�,���/��*B.��sM�gvQ��^I��DR�g�bġ�3�����@���ߢ�o��gl�)S����^(�h���:�b�Ɖ��@�C����+Q�\�n�녙蚭��\�I`[ѓ� E������<�� ��� A�~}[��.����L�)���X��/!��6�K��P��k��	���G���!��^�����m�F�8׼��mͮ��a��>�)S_�
L��Kw^O�=�-v7;f(�T��Zv�J���s����H%25�z���lx�y��s�{��D���@�L1��Ԙgj�=���bnϺ!`���Yw^��T�O����)��Ԕ�b��h��"r�-���@lL�5�A���AoC6]t�K����I����G�Sύ!=rr��/��������/W2K��o
�-h��T���/��\�$��"���K�]ޫQ#��KB߻4��7��'zɱ�p`��@��e�C��AWΩ�$���ڊR��u����f����ϱ��jlS�w�Z8�]�BSR�۸γ{�͙J9�񄫵���t�:�ҺP�����I�;re�f�8/�Y,f�H�w��pr�u�dO��E+�3xCe��@��"�;��M!-�^4�ܫ%^Kl1;~O�N�1[
���E��	��k��7�1�3��Ȭ����Xn���oP(=u��luq�Lgn����KkV`v��)���x^��n���4G��`"W�����&���}M�x�+U/ J�ƅ8�4��s����=ͫTw�[��-���-�Y���E?�pץ�?���[����7���K�_vp�1P��(Z��	M���g���փ���ѻ	���	Z��g4�ȦP��8��q��M=x�b��0���e����t&5���?������X\Ҳ�-���z��8����n�C�8�(.���X?w� $:"���_��%/�f��{h��G���m����*wX!6f l%u��W!A��4�f����7��WC*���XF�eg҉r{x.��oT��@��Gr�b�0�Ij������1?!��ʓ��k2�e�B	��j��6`�(�j�7����O�����a��*�9v2�R��1 �_����ֵ�����7	߲^hH�|�َi��=7�>c�|42q^��]a/�k�3~��l���^��c�Ƣh�F��%����7�1I�BO����
��t�fy�ַ�E~�I}���жs~�1'��T��"QSOV����U�O�a����#�z���0a?��OQ�%>=�o�/�F/��@�"3N��c�G��d�ʲ�!�HEt�n��Ԝ�ƾ������c�8��&h�ݺ�l,���5
?��=��(O K����+.�V���^V�.�nI	���'�?��(O��=�=�qǸ쎃�q�t����M7�<c�ݚ3I����'��4��((�a�����2��<��:"_�E���,�.�Fa[%ș_�([ж[j��-/R��^�LJ���гV�<X��Gs$�dY�q���zq���_TA���B�7f�r�mN���:Y��q(Wj5x[1��U!�F�|k;��ԁX4���6xM~�u�� �V;7��E�Z�	���T���~dk�J�� yΑ���	'R��J<���D��E^l$���UdB��HM� �Ύ����n�� ��}Mk�]�= ��}�/�J��ڢL�Z�.�iA9${ӈN���3�ֿ
��%�
�[G-�)����+�����f��ح��i(�g�՛l�T'�Ps�V���罒(��ʪr�=�'��9��2|̗�� �M�ɑ/GO�55���=k�Hh]��b��~��w5�i�	���"d��ԡ��⏳b�p	:G�FV���|�"�I6!,X���/MƦb8O��^�� ���1GU��1�uY�=�b��1�Ȏ���6E�L�������q
Z.Pi�{3ܤ�PQ��7kN�F�0�|����gw!N�*��7,�W%��}V 2�)��Ū�J;��b�P|�#>P	:�4�K\f�4�ө��^�Mԑ��,��5������]V � H�_��|R:�dv�x���+}e>h���^hVH��o[�vK�.����M.h��Ju�]R��.5�D��{� �����`*����&ʆ�jp���;�aS�e�ZF�1X��˂ 2���
C�%�2�+'ӖF���eF���&�	�ח1kA�|X��B�S�q���}]1m��`R�&�c Y~��S���W���O������!�4 ���R��\��
ĸ�}��?�)�-}�\�Rq�w6r���@,��,~6�z"���a׽���E� �]�g��{�%Yq����EO�����U�%72gE�ZVUv	ؘ]H�1����� ���-*t-��k,�������ܹ=M�`��%��T�oPb����P �����l]�T��k��1RN,M)0�b�j�=�>B�s�ˑ� �|4�C$*��k�,�����+<)2C�=��Ƅ0� V���������=#Q'���h����U��{9�!��.�+|>7��_s�)�Bi�gPlE�L�$�����|!���/{UG��R��P7B��ovYa�=�i���~g�7�H�	f�2z���d�ŀl)��42�86�rrѫ��HZ�y̐�l$XH}��/^.m��r"���Jd��\��f����^��S���� �0zE����1>ݛII�yU�U�M�C�û�$&�"�!	X����*H�Z�d���w4���T����1�r��uZ�;����(���;ؗL~���ia�"��9mh�5��8v���03p�Ph߸���T�l�����X���D|0����i��tGE�t '-䉍���Y�K��������z�1]���l�/��)�  L����e(n��3_VQ%`��z�d���"��S6���W�È��ň��B�mQ`v�rt�*X���77�~�hX!���o=
U�E�o�S�Oj7�tO��#Y���A�i,i�}���!�����۸����-n�-sv>��	dhҁ_���nKĿ���':��V:"4��g�e'!�:��>|�`eu
uq>�y������x<�k��vWi> �3��f0)��1���'B�M93e�؍���S�=�s��NP�W�	���Iw�"���ČoH�N�u��$g^5#Wo,�;�Y�W�d�T�&!�&U��o�7����i�y�WK�
E=�ʹV�����)�c��T�5��M����>ѕ�K�ɂ3�`R��x	�/�@c�_�lۦyՈi�+'��
�N-ջq
���;DhIέ�󤍖��3�U1uW��&kJ��PTԏ�L��ӯ�K���l?ؔ׸����h�O�:��p]��z�7ޫ�Im��J3$�N����M3ϱ���a*��:��\%�O,Dg��Ԟ����Q�%�Vq-�^,[��tD�r�?1U�l�P$6$6΃��u����*���ߤ�t�+��9�.���2���:���<�*��YT�[��%O7�[U$?=�-Q�����++��=t��Q��t�=x&�=���݀�?U�b��*����<X���Lh��ϕ�G��I94*��� S-�*p�UUQ��	yT�-@�;ٻ}��7XzH'rB�L7��FI�[�A��m�����}n�m��ݻ�/�g����1ѥ(k���j!��(�7>M��r"�y�ۅ�-�L�C�t��= ��K1�D=DW��omk'�jaq���9�Z\ n��;y�����$�;Z庢�h��\�Li��Wio���d/���Լh��U���`6��'��C?��1�c��R�L��vț���+��s��Ü���Z�G�d�� ��s���w�%ѹ��k�>e���M��d��Y�~�!������=7�C�-&᧤���cĜ�����l�oq��/5����a&U\�.G����v-��x�o�o;�[�e��0;���#���