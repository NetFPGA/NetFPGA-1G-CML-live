XlxV64EB    20e1     b40k�s��̸I6��M|�����p�*P�\�~�$�+;�_^רL��,����$������}�C+}=�Q0_M�'VQX���4M��E��Á�-���2��~ӂ
r[�bb4���R7�C�q�k�$�ї
����1�9�m/����"ב�@����"O~�xN�ܫR$���!�r-$��~��9���#�����Av�l�����J9��\�B�i�`���,V3��k������w�K��%x}�aj✕��U�]�@�ۛ�:=�JR�AA�3���u+p�VT2�����c׆\s!��D��#��>>Ķ����y���_O�w7��]��xb ��p^l�A��FJ~��SH؁ϧ�{n�����/�.[$ ��wA$��;�[N���Ah�d$��A���+��:�`��F�FQO��jǕ9�1B4��	nƊ=�����J,(K��Ԉ�(���'��L�D�����>g��0���ˎ$�2��G:]�o�5I��I�Ga3e�8c'[�¤�Iv��f�|gb���&i�LGL�Y( I\w:b��4����fP���H��c��Θ��}��/gD8�"ZB����r��إ�>�廊I����#�%�[�S��6m�����P9��e���L�g��m�U���]����u�{��^���$�CW���k�.��)�봮�:�Fh˼ĕ��ي䆢T����u*W���9�Ԙ��q�D��QP!�B;/��Z9��_ګ����(�����;�3�k�ރ�`����tQ���eF���S�	- �C	o[�MVEh/k�	���;�'畍�<���W�V���ޒ"#P���ё���+'K����=�ZP��<K� J���l��A���2na��w/V	��n�o�e�9؏K}���E�^�1����+ǲfz��j��3'y�zւ�e���<`<I��a���a����0w]��n��i�m1b�_$;��N���x��)��'�i�F�<8�����l�(��i%�!�؀z�q0�@ӯ����<�=��q��s�w�N�ğ%�lF������_������S/���c&�FzZVK�H���G��.iW���G�����<|0ǖ���8���*�3���qᨡ�L	>>
϶�ݝy��47�#�p�q.*N������WYMY�D���B�c�����@8��*
�R��-�j X�L�[J�Gs��%.q:NF���f�&1����ȷ9J��si:��;_�>�FqA��Q���ƺH��N�(�y��Dڮ�C��ۮP'�;����̷jb��mE���D�96-��T��1H*,PB��O�P9�B��#4�b�X�^1��SNi�RQ#��ߝI4���.��`��?_����5_���ӝzt��FyK�E�6ԣ�9���H��}D�q��u��]�@kE�«����!��_�� �~I�C}��F�zk>�!�/
-��-�?��q�2�yY��s#V�M�RM��(s�_nAM����x�˲`���/���?��2�'����3���W�K���\EF�g)�D�G�:O�"��ј����kO8����4iT�2�H�H��@��S-����!��T)��u�v�3��3���9�py�XWP�����܍�C]1я�P{TkjI�I����a�#�{6���[
C)��y?C�+�����]c� {7f��LVtB�C�~N����T�_[��a�l�2�)�L�χ:|��5cpG�f��Nt
�2�������J��p?�sɠ}�}cu�[�?�AJ��l��)����ri�Q���c<��W�*�<;gT�^ӆ��d�k^�x
ѕ��^�70���l��0%�"�+�\��4����r�q������Z�������`�ՋS��|ڒ\�xț�Y\�^�;Ez/	 n����E��p|?+ \fy�_A�������6l���^@��]��0�6P�"wk��Ù����#a�c���x(���'���E?�����iZ`.3�)���=�ٙ�u%�Hɕ�xa�p)��#�{��s�q\?b��d��}�&�v�ߥ!#캨�d�PU���0����.�0��HN�0)N3��h'=�
�{�Ru|J[|�"&�a5�����y?�6Yu]"����9�(�|*�6ِ��\)��������&�=��ni��g�O��<+;�3��\0~Wռ՟����ydv�c���;����� 
�0G�to�\�S���\$����M��	�hN���2�f��Ҝ�L��w�����9�4����F�epk���,5`��\gOq��x1M�o�/۪����9י�᱓�pN�9�Swάd���E�+����[3 �%_��a�j��Ui��}MX��L*�?�ɐ��g�T�z���NeC�S�KsXj�A��<���r�GeV���'ĿK���j@��گ�-]�/��������٨[)QJy�$����:@ǅ���O�Mq&�J�9��8��ᆴ�r#ԊK���y���%�EX�;�I�mc��I��iݿ��[��k���W
a�ϲ[3wk�O���KJ7@��sP�Va�=��ﬨj�j:zt�K��xaǞkφ2I޻,	Hŗ\AT�!X��?�W���\eD��Z�>B9��ъDiF�l<�9ZM�D/o�e�<ߠ�S�ػ�#����ǥܓG-Y��yڐ��)�߳���	����n�@Ʉ3�y�A�y*��)#r���'���b�7�M���h�`R���7�/yo���_r�	�v��@��G$ʚ͕��Er_$�@�볕��Z��Ed�����2