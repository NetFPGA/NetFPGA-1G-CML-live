XlxV64EB    1b5b     9e0RA�H���jF�9�Ih�6T����q�����+C����blo�J�쏲n���GT�_�/�Zʬ�)����va
e����V�@��&?0I&N��� ޠ���3N�]�3��<� �N9j�oQ{���@ɺ�خ�i$�Ф�,��v��N�Ǩ��)s�~�ш=�<x��xo��T�q�d�n՚C����bD���0��nc
�ڤ���b�a�:�b۫2��l�.��AA�G&ȹ�|�S"��$�o�W���C7pm��E�a�&�s�uhgF�Y�e����'u-~ڈ��W(���x4��s�S+S�ۈq7^W�~Kaee�A����lj!���@&ҋ���σ�*�'|_����Q���]s��<�Ǹ)�?]�H�R`}i��� ���+�9��?"]�pV�<�>H����FN�<�7�m@�b;��τi*��yj!*�ᩭ��VڽH}%g1$2u�9mm��O-qY��J�RDw`*=�w��V��i]���T6��|��uO���
�;��+J���
Z ����,'ł�Ca�;�k��
d+�lr�1��z����M�GE�X�2�g�p�2C0z'M�r���.�4=��M(�
�G�4�t/�B{-��W�k�����$^��>O��^�ݙ�p*��a>�r� ��nW	I\�*���>�3���x���.]��u�1���#Zb���&&� �a��?7��%������� O�fQ@��\#�1��V"�0C9B��ˇ�*Bơv�Ůs"��e��9��A�r�Ch���E�ɣ��H�_�*h�,�]��7�%���٤�:�`bo?�3���ܞ?�;��R.��ʟ���������I���Zփ��P�^���I�ɟ!� ����g�|�2��pzI�����{3l|NjǯA.y���SD,މ��
ٝY��F�<�!��~�ONФ6�nh����W�P{��I0��6�ۃj��D�oI�­;�Iq�L���ȭ��H,��~��Jb+>U3m�=]��]'SS�O$C��֖�k/]gYI}m&h2�M��(~~PO�?T5����Q{����8DE�G����{`2+B`���΀��UL�} E]I
�|QFq�{�J��-�!z��}$�G%��1Z����ҰC(,�<�9��)�J`4wM��'� �� f_�-�)�|�M� $�ɛ�	v�b+��R��:l�.�41"kMb�bA�����sAil9�gD-46ʰx�w��������B�%��ިy�e���ֈ���a�m���`�-��Z�;���F(����֚X|���~�:�"�E��ˡ�&�3����~<Y��̨��}*5z��H�*,�!	�%WȌ>���.�V��j���j3vQ�]FOl�d�+��&�a�c��8�uc
��7?�L2��so�l�Q�Zi��hЭ�+�Q�x-�e�A������Cx"�h���8 ����w=pp�ts�D4 j�g�՜R��GCs#�
?�w�QQ�L~��H�	I��FM~����F�G���1�^ڍd�����y<��a�9���l6]��������K`K��57��i׷���cIP�^��l�Ov��l�kZ�g7���6���_P�̽�;��?�ZrKvp�iv���{�F�b6ȩRj�Rݡ�y��Ei��/H�=�d���N̔�k�%a�r���[.�
������m�(v%�ߥ6����{��R$.��:�+��}>�j�]�,6-��xy	R�����8�/Y���N��@����6�?�^X����&G:����)r�T3mǠ�*��Ű�Z�H�n�y�K/�О]�2n�ĭ���`-��&��F��ăL��cLyT*�ܼ���_�/h�������m�2_hx�~R��/2�,�+an�Bg�bC:e q�K�͍o��{E��ڊ3+yH�1�6&��j�
hK����m3�.���G^M>�H�~D� @���I�D+sEO"rU^i���<5e`nAx�FtKKD�	S�:�l|��+b������s]c��N�cjH�$l�c܀���jɻ`d*���l,�:��ɾ��'����V��!��+�A-�M�n���Zn!j|=E5��s/�\|��__S��J$�יS@�Z��ă_������� �m8>74T���W]�?��=Q�s�٠a�0�{��eY������Q��F�5��Ϛ�A$�|y'�G�j�l�u�0���l��OE�3���@����׉��
��Nu�۲Zfp4'�O����eB�V`�QĎ.�.$���z���|n�6�	4����;�Um
�j�a���q��$�Sh����]��mOP�ͩ�7ZH�H�\����]��Ֆ�;i���X̿��*�Q!5П��0cu��t�������5A���Q) �g;ߣs��(�Y㮏�x�zj�d����@Z���}�a?��>���
���2��)}:S!��|�eŵ�2�i��r