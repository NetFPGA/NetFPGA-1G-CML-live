XlxV64EB    2459     b40�3��9�� ���������zДGQ��A�Ѕ�B��A���H0�'۴�5W���=��oϙw�K��!C�:������0���m��
'K�|��K��D���[��Ŧؾ��$�~�/4t�j�x�k�N��{��"�$IVgT�u(yJ�d��2m2�@�2E�C�g�_E���<�t�tZ Y���E���9誳�(
���4��8\�X�9�Q��H���"Y�+}�c����N�!s!���a���1�T�:��ݓ=(#6��Z��d]F���P�kvTp�)}����k̴dq���\�䱇I��q�)e�َ��|�!��&׵�&j&���'u|�4��a��Ah�S���:����"ІJC�7/e���G�
���hū���E�5d��%���ϭJ�`�n��g��u�(@����zwMc7�Uf~���*W���o�� ��B��g�f
�-�����w�KGk`r����9��9G�}� �F�;�g��|�Jnꠖ��h�?�6Pwa@2+@���k��i����a0G��T~�EL,�}�M���[���gg���-�D	͑�ΆH]c�(7��'�#���ڲ��.����2*�n�H:t��aL�}�6��?2�����?�iq���G�B/�K�8�X|Z
�m�t��<�h�z�h�q�f ���!fш��t� Sw�w2_R���Gu��h���oT	�&1x&�8����3�V?�h���"�hv�l8>y��iv�!^xؘ�x��9��kd:���m�r�'3��UB���2���	�5���t`MM�S���?��|�������L�2����X#L?�+i�����T�B
��=ͼ�u��/ ������Ͱ���~������2z��ݱh�i��?�2��t�*ЩQ���xuirz��Q��$f�Ԯδ������nr�Ty�Q�{ߖOg�j*���*�o��{ȼ��4�g��O���,���ɫTL�/0��i�]����N�
�{!��a��LfE���C��m`�	�[M�Ir��F���r���<�,
�S��bu땍B*`��ɾ�Hjߪ����1��91�7���֮���SW�4(�槂8N��Qg��_����I�mxD�����2V���� '�O��'o�Uo:[�+��c2����rZT(�DE"�tD|�����-�X�Y����H*]��2�n�T5go�z��ʨ'|�~b�jD���bB�-e�.��N�
� �iM�� y�����0Π�ˮu�A��q��Ֆ�n�U6���/��\О^%K0��_�si���X"j!�t�]_����`�uo��ˮS��#p3>�8���y3�%��*�J_���RG!�V���㫵i��M�~m4� �2&��΋�X���v��`��U+K�����h�$�	黅_�������.�0���_}W八��6CIO-�a��N=�l�-f0Z��OdS�SaJJR�a�&}f����Ӆ����������nr��)����������"�FQP!�&��Cϡ�suj��F�j�O�0�����ז�*S�1mþW�4Y��i?a�����Պ���'k_�U;`�Z�qV)\����!3';�� ��1����f�YM}�<$�!JI?��|����+�o����ؚ/V�H�����'��н�ԆFw���w8簜mP�:�j;���?����x��?�=��zX�k�F_ΗO�T*�?��Ud~���]�O\s���:�A�&Gbҁ�h"�5��0g���Z��M9���K1� -���Z&r��(��F-4y7B�]o��;�_Ӆ}ݒ���n�w��	��k�T��W<��<x�F{{�>c��v�<l�T(�Q�	�S%�J]I��>��ߌ����9I�-m�C<�I�+.ǰ&�}E#M���rޭ2ַw�G&.0��<��Qr�U �!��� �04.i;_q��g(�&@��onC���)g�oS���A�Ab� ���R+�!㈞�`zZ(����3�ͶPp���4������J���s0��e9;`�-U4���Nt)��u�S������.b�$&����r�c�P�s���4����W
�����Z`�7QL-�{�O&՛��&b�5�Fs�Ĳ�E8���M��{�^�<��c	�I�3W$��H�~ �8϶c��Z��T��*z}X{��La�'~��Ư��/��MV��:l8����4�xR!U
Y���w$ʴg(�V�͝�f�i{ ���q����B��gB�S���To�ю�~�B7�vk�+?�x�A`��]U�M�������[Vx����>)��0�����Z�t�W��y��"�ȩj>�Z����@n���s�z���^�4�i6+�;�m���8$�!Q��=�zD��M�(���$c�h�f�S�d���5D�ݻQ=l�)��Bo�������/�!r��*��.�G��u��3�6��
��i/F��� �_GK�Kw�����E{ݩ�1ZS�	�%���h��CW��e��������'f�P]F�AGf�(:�dqĕ�����m����][�S��`�r��ے^꫹�bj�7��Er�c�����15�w��}�	xŅ��s�+k[�qݘ���ă��: |],W�zp:�~~�rm�(��0�[e������C�"˸F�6����a�M�8�N{� ��tt���Ը�,3�y=�H�p4t/ԇ���c��>���|�+�.�&A)��� �c���@���}w��1���[�\�k�I��-T�`t��xX�L�f����Z3���cn*