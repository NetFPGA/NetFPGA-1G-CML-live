XlxV64EB    55ea    12f0
0;:���f_)l�dzN.+�'���Sw�SŦ������rK�&�b����L�t�V��$�6J�繑;sχ��������n=e>T���5$e��=y�w��*�D��DO��o��'���T���4�87	�4ňh�!�\59؟q%R�|M�q���%�c��/C#'�e�;A:1��H��y��IW��E����A�=���ϯ�B2�Jm�2�o����$>ㆥ��� �X7t��0����QV!I
m|���+��wz� ����Kwr0+4��T$y��PEU�z]�m���mQ�$����(s��,黧|7 7�,����Zś��~<�{R����g+o�l]�/��и� g��;�&�C�������o�u�ju��2�I�0oE}�n�k]hԲG�P�(ef��'uM]h��r�t\,��1d����L�;c��+&��-����>;%������DGY ����� �7��I���a��Zk^m�봊��E_�i-����k럗5��1���Z��%�����Y+j;�j��KH(W22"�����:%�T����_u��:��C�J �~���:�s�HN�K֕-��L��v�+�u�o��*�.�X��|H���Vh�C#�s�pЊ��M�Uߦ.:*L��w�`j����;CXBiAK�ٙ����<������鳫^m�7�����>N�D |i��Z�����>�7�������,�H����Jj�o���N%�([���Z�# ��u\oqBeY�+�a�c��D,�+L�q�v�)gZ�5���F�1ic:����6`�.��}�jOh8�y-ta���P�Qx�ƭ���x���L�ؘ��)$Wzzky��8\��c�=�oKP{�29�u#̤�2�1sԠ���w�;'~΄��9O��8�X�jic؟:��,�؇;}�F�\ů�&��H-�+�Zn.9����1����r�Ȯٟ~��^T�7J�5�������	$��;n���4릂�@F�>�h�#Ѱ
G�9�����n�N�ɶ�q���O��R �ZUJs�������a?%��0�ZGl�BR`R8y�4ь���76@���x4���ޭxl���e0�. �
c��˕s�Ǜ�����[zO��P���2�8#|�(� u����'8҅#�iE�!��*Y	dϜ/C�cכ��E���d0�&���&lT��*][�H)��+��c��ppA�6�$���V��qjRJ[w����|�Ȝ�!��i���#ֳ��4�;r|	,�lޤҦ�W�c�,U��*�6�sp9�4��?�t%�!ui��˺�z`L��q��E�? ƪQ�)R���b�^ǮGj<���g���>SK�TL Ϯ7���>w�1a�߃���,͡ߌ��}��<�$��~�
�J�e�ʳ;ܑ_��ط�O�*��'��ڐ'�� rձ5����×nX���W��(c���b�x�d��AV�b��`Rܴ��F._]�|��ѬLӕf�J�p)�Y�ON\7�@� ;z��4nlkʔ����0��6���',y{;�d�$�>��O
�]�i�:���D;5�f2�cU��n���S�����l�U�����{4Vo�|�wZ�����F�u��z:۠�#L���[���Gr�v�5_�G0�͒ǽ?�#i\O�t�_����Vvu�S����
Kq�:Nw�D��3�ń2W}��Q\�/��J`����D9�T��.;d��&?�*�>�\,�8prNʀ�_+>EaR�����+�f�"��$�b-ụ̏����I�Mw�^+@�ԉ�׼�!�:����𧲔��#�!�/+��)�S%W���ծ����Ǧ����|���^ҿ�M��9��������e+��E�<���T왟[`��n�i�W�^�1�1}�r�Q&T��tre��2�7���>�_�K�ʨ����0�V�Q�hq��0D����� ������>�0����WEt�l����	m
K�?_f*�_>�<g��)\��al��2���k��z4��}Dv���p��Mf�۠D�Nq���`e���R�էn/��0N�58�� #T�	QQgY7.��$�6Ύ��[ѫŅo��x�-�%��N���9t�_�yx 8�wr=:�"Ӽ:E��;����*�p�ȹ�C��Ԡ�����KK���W�R��� �D���X�> �+�_�t���78��6��,JZ\
w4��J�R�ܐ�̖\��>��X
+ޙj�0scc5�s�u��Y���~��7�?����T��1��K�-�%gº-�mu��N�֟*��A#:K�'� ����NR�����qw����zdx��c��kΐ�&��[� &�"�ːչ@M'eۧ����ܽ���Y��?����)b�OW�V���#|�b`"��~��+f��hJ�Q3�!n��
g�c���n~K�M`��S.A5�B�Ac<^�] ^{�>_�p-7COrI��|���eO�O� ����9,"��czj1��|n�/"�e?z�����"z���1�UF�<��U���x.�{�k�pF�%�ذ�m䣮ݏ�N�������Kms�T*�(*=�v���Y�T�.�4��E�w4��թ�T{�uS��K3���s�3�X�+���z �IM��%8$�Qu4�-5�
�'� GK�\ş4�ΛBPU���0�����:ٶ�����(��j������'�.GO��މ���i�a�=p����#)v	YMfE�.����٧1w'A�e.��]�M��綢�{\8���'�5V�}¤M�b��~����OiK�m3���X��S^���H $V�/�ꪒ䅆�rؖ�c�[}�4
s�:@&�� e��A��둖+!�ɾg;�y�.��tw�6J[4��'�x��
�u�O�8}~��}�iw�!���g2����+��ϭ�,i��.��<x]��X�`�����"6������me����v��;LlA��_����4����Jt�����hѭ9��+f����`�S!���_�V��\�X��Z	�B��q:�\F�'�fs!a)�
K��!�'ѻ�&{	
�F%;V.-��&�=q��!���Ѷtb(��:j�^��#��X���"N@e�zce�b����d�՛s��2�3�otZw����>G��F#�����9���_I�y�?�w|@�V`�_�'5Y���o~f� ���܁��;d����v����z8��>��ڨ�?ƌ��i�}�����R2����X��"^����"3���M��Ŀ�}o�r1�j����Q.'xJE�A$��&P��3����י�W�V�A@�,�FU���������3_����*u����:j�����
+� K�[��1�h���}{���9y�J���yC@� wh/�߀�J�N�a]0�y���ܖ�@�9ٚ�p':Tbs���J4޲p:�l|���E��l�T�&wY�1��>��s�)D���y5V���!y��D�|It�f��e�0l�#{�*�L�a�*N,�.�]���tm9�8$��23�or��"S�;��;ZM�(����ꋟXj�:rG<L�tD�c��ȁ��W�Qד�
�|�ޢ�F�t���͘AJ��r5@�jM��}>���:��k���Pi�l��M���$fu���v���MĊ`��͹=��Gm��=��|�]eb=�}������2����#?��?BF��*����Q٢��r�_�'��e�Z7)Ѻ|jg�]�lϟ�"��l�Ϊ�{�[��8v���U���(*���k��N����i��t��^m��Q���?���B�D���㢉��e�r9d�<cq�+ME�@*���r�,Q� �C�}���09Q��yb	�XM������q�6�"ɯ�WI1�E�D�tT8LG�3h��߆��]l�P�2����+�{��K����9��O���뽐WD��x����Bķ.Ҏ���|c���=�~���N������E�����AiŲ�U���{�.w���u�󤬱A]�qX�/Iv�)�N�ck�4�<ذ";��L�^BA�~��K�\�-{P�˽'4�M�(�ɤ�JHˈ����D9Fw��h���ߊ��!� ��	����S�g���z(�Ny��U�T�������Av%�7�=gZu��o"�(UI�_J:�D�<Z�w�KR�QSC�>�rOm����p�(��yD0�x��2ﯢm�w�Hs*&�*��.7Bq]�ea��)\mW��C����Vz$�6e�����H~0?E	�lBtI��;"�4B;����GO��a �4Ӹw�B�G�6U+����^����2A5�h��eWǈcc�n92��H�q$�<�u��84&��,�<e�OEŝ/E�p9V�О*��u�Iv��A�%��u�!8�����tb�ݓz�Y�k-_W+b^$�� �Q3?er-��-��Ԃ ���w)Q�`8sqpȶ�!���4ϾkPQY0�i�ǚ����3FM�!�o�;���p^��nޓL�Ǖ��O0��̆��)I@ڮ8-��������t�~Y����mzV{"�:���2U��7��oޤ�����D�C��3HE��V�O7��t�Vn�p�8Ș������M,i$�<Wh{�]�m�Pcq<N��z����"�8���-��'`��.u�ɕh�	 ����MJ}]�6����m�q��q�w�\���w@��F9d����t6�o�