XlxV64EB    1b83     9c05��R�=H���@���:���9`�=	�hzqb�����	Y�hf�T����Ym�=�ճ>�\��>5jB�F�g3(I��+h�Z3u	��:�E��̗6�s �Tf��YmZ>�tpw�������)%�C�D%U	ߍ�g�zX��A-�oqsR�F��	��'����*�9�柏�g�{j^K@�=DM�\GT��kj|���<+K�DY(-��#��)g6*A���H��7��V�D��J�� ș��Eg,H���,��{T�b��j��8,e%dx۪kW�����O��@�2��u�4���_�YOJm�+�4=����֓���/r� Iei�*.*��;�)]���+ ����\e��*8��e�#]���B	y��6�;yIY��38q�O�0X���`P?���P�<g}v?'�d���xPҕ2p�LX�Z��2x�����{W� ����!n���}���O�\�E���$��X��
�Հ��
��d�SA�hHh��p� ���9�+�"��3 �����n~`G@��=�BF��e9�O�c7����,֟�ig����+;т��8�)k���o*���=?��DD	<c�f�HA	;|	���+H8��ᣄQa/F�����c�"X�(M0���3�f[y�ԍ@޷�7����]nK�Xԩx���T5�W�5�j����A��8TE�s٧�9D�+:�U`6��"8��z�5
iF�6��Y�t)!X����m��32�1�J#&��B��M.��N�x��M�.�5�+͓�.P�C�@aQ~��:d:��sķ�W_7�C����#Io��%�����^I�A��xM�H��kU�H����S)�k�EszJ�-H��^x�� °�Ȉ[�:�t4�'���8�����Փ\B4�qS�He$��O�|��Ș�W�n���oq�����ѷ����{b����QN/��D�Svw��;��2�J�<�����p�j���*Z}\E�������IsL��>IXH������L�Æf��Б�ɫ����ʺ�@�����fL����t9y?�A��u8���cT!,���㩸Ԇ�E�8f��BMi��\����I�iTaݜKy�wudRz�?/�4��tq�α�>-��KT�bc#c�G��b���\b?�&���Ɍwn���Kە���WG�����c^Eн����u�N�z%I�U�}�����O��=
U��R�ؠ:�����C� �f�p4�V���~ܰkD%f�#�x��L���Dv�d�jxJ���K�fK��j��e��d{z��dy�&�BDN�xH���P���J��7��&N��;��;��Kk:D���p�Y ���>�-U���bBB@r�y�և쒣�oڷE@�YG4I�c���� oMɕ��FQUtS՟�s&k��u�쎼�H��oI�A�4��ϣ-g
��M������&�|���P�ȕƶ�a����a���S
��9p���x��/��'&ӐWIΧ+ �/�R��� 2���t���Psܲ�0s@n2�L ���@���}�Dm]�9ڞH9G+Lr%;��_�ƌ:$R�@eK���l�Jq��7!�N�&���MF�/�]���.	�NF�"Uǻh�#��q�T-������P��G=6��j�k{�p�8pZ|��fL���m���5x�c�)�Tڲd�zM7�>E�C����L ��oB�da-\�C���]MJ�1��0�	�R��'�����u�k��A�7�O���[/q|���3+��'F���F��Ur�-�r���E�31�	��a��e#������q�I�Qܮ"�*e.�*߳���gf��qi�R�����)�A`��dIj2�ѐ�a�ԍ�=v��|kU��$.��|L^asl�����YcU�hvSn�D]��z�֗�F�͆���}�/�5y/���
}�쩜5���,)�>�W������O��0��x�	?g�R��K(�}����ʀ�����t��͚PQq�۱����6� F���������W�L��5��o���~M���#�ɼ�eQ@�PT-���3y�.jԣCY��S�2��+s}�9��r��9�K�\s�K�yc��&
���s#��-�g�{/D�Sw���v�]t����Dd�������HAJ��*�!j�m�w>�O�e����1�h��S�9ɉ�z8��7R)OQ��?Ib�ń�"^��,ЖF��6�W]/�}�k���B�J�\f6Kg>[�"D2Y��t^�)H�f^9ёm3�ɱ�/�V��w��DLWc�?�����5�m��u�L1�X�OsL��~2	�����ꪷxҧ�Ts�C�P������=M״��)�C���K�:�]wx��vf�J���?ETB_wi��dB�'Bt���Z�yG8���]hM--L�0���f��RH�� ,O��~�zP7�x�࢐��7(�*��[��F