XlxV64EB    fa00    2eb0�
��q��S�du_�#F�l�䑅63:\u���j��/�n*�܊��O3��U��Z��YEn�I!cC��%���[�4�l����M��*��=(Dqưo�G`9X���5���t~�q�e�~t�#��G��%��Q�P��<�b����AF�S����5ym�˴��ע����H��dË��B�
�8�,m�G`��>2��������� Yp�cz�~�*L�X���3;_JCL�j���ْw�t�|���v��>$7�x�_ټ+u.Ac�K0���܄K2h�q�ZbN��{5eέ��ֳ�0�b�e2hm%&3bq�[�̭��/�>���"�Y�dwz��C��{X2�6�ˮ	��V4��Y/EzWϩ��>�Wbҽ'�����"�"�G�f�����dwz�C3������b�I�p^K�m�T�9z�����;$�����l���b�I�B�xx��V��"~k5~H�� �Q�c\V�mXS�a�q�݉P�Yw�w6E2�8��rc �%���U������c����ؿ���:ԮeH=��-e������z-;6�:g�B�ޤ���)�����KL�E���̪!���Ħ����")5��/k�7��}�����vwy�oZ����ސ��Tj�Y'�x�O�|H�������!�%3Vxܣ6`�[�6���#7�������t7�2����q�rB̧a� ����{03;�|a��*�v>8��j|ƥ����5��ev�=�>H:�_��P9l�9s��E;�3e��F]�������41P�e����\WF�!vx���.qeӅz�y�7����t�V���Q�ۚ7ūּCe�[6i!����쩞��'�����|�)qG�~0��GmƆG5	�~(�ZF˼�Q��W�V��-�w�DJ�%�����M�j
U����� ��W߭'�V8��d�Ԁ����j���-�F�2ߺ��S��򪻽�9�uﴧ�y6R��Y�|����R���.�t��	.��-�)�B�����U�B�EW����	.WM��٫u�w�u!�ro�s���	��jS��?/5*���BR`�����zXv�����jN�ϓ�w4} ��&5"qZ3����CR3kѝjP-/6�[��p�M�&�yM�f��r@��K�4�=���9Ta��Y�3��}
�p���_l�@4W�{��`�$���y�-��y�*����#o�Ţ?�O�1���������]]9RPR��+����z�(�8X�1�;X��'���'�$m��}��*h�v�(d�#�ќ����KW�T���͖�ƧX𸈖����&^�p��@f�]��>M��J7�C��-�Crt���zgx�^�ۿ ����PT|�Xn9�@)\� f�8��Gu�֩�+?m@T���e}1�_K�:s?��*p�r����=�\3�������ŕ=��\� (��sp��t�!�Ś�f�[z�p�k�T~;��l4Ku������j�x�Aoܸ�b��0�d�.��[Z��V{�	8݊�(����I����d��^����K��[�[d�@ a�r/J�n�]�����Vv�q���U_�72{GR�M{O����!/E#2BPǹ�MG����� �ٙ'�i�W���,4��������E/�<@��,�t��y�(�,��X�-�<ݢr�)Ǿ��P���^�k�\���$z�޲TuWwD���	��H) ,����o)rLV�}�n=γU=��*}̱�$0i�+�4���Bs���9CЬ:vt�W�T�9Iⶩ8�?H*��BK�Va��x@�[ŪW�5M��'�� X0�<0  QO�Tj�<&��e"a�TӠ��yrv��g
��՗�a����<�
ϭ�R�(kx_�s?qݴ��?F"6�í{R�&CjnN������㊖j�咙P�q4��Y��{#���#AT�����M��|+D�i��m�)��`.�[�Ao;�����L�>��ߔ��.:5�nG��5�L��"'�%�e� b(S�l���6Mt �]H�#����O0�����oW�3��=���wg�$�����}��"
����ب
�<�����5	�h���4�� �uCN�iVj��%b��42��ܩ�C%D�m��������U��E:���4�1����r�s�v�𠔞,(�c2��7I���VO&��m&q����/q>�%<5;�+8N���'{wrU�05A9�U�!�� ��)R�r�f��VL���e��g��ޯ��W�gv/J��@�}���T��a��l܁����9�lX5�)�EQ*��N�=s.\���;پ�_��~��0��:�L8�H�U��e����dH>`E�&~�� @~�΍���N�-��b��:�mX�i%�Ay�$pm7��%�г6港��Jj� �aXI`��S ��W¼��G���Y�y~�֦��[eձ�9�?��/��!�TM�L���NΒ��@v��3OJ�)�TbGTe�T�t��=�/6㵕;�i�uR��㖩o��&2MM|�<G�����B����Ke��J�;�<�t�2�g|��ɾ�]��vҗ`�a���7��b�7�҅-kϭ��O:_,HJ���ͷp���_�e��X�`!��2~рVZOC�k�{�J���s��j��r��\[ց
Xl��9f�8Z�O�R��&\?G��Jۓ�M���=��W<Z�ȫ�L! ܥH�@��-�ZL�B�I�/��xe"▖9����B]�@1���u����Π�7[q�vݞ?M����f	�a�g���F�
/w�C=��Pɿeљ*�u`�c��`��?r�=CCC�4
H�9�MxEg����3$�f7�6]�k�ͱ!I51₁UFfA��r�j���w'0}�r��Fƣ�lq����ȘA����V�V@T���D@G�%&�
u�T������y� t<��ly�O�>�MW[5"��λ�%r=ӻ�ln���_���>��QB���p%��>��!��4��<^�_�G�R�߰`��W���p�c!��]�`k����ص��c�%�T[��x������ܝ *c���r����
��Y�~r_1}p����4i.;�qI&�l.#�;7�d.��4��./]��Q���U<Θ���]&��6RO{�k��&tz�1�uğ�sD$��g-��S�0�XOp�q7x7�����vO�!a+�ɢ9F�D�V
�>
�R}T��S,�ޔn��������I�-��+�Q}s�o��Z!��Q�{�+�׀Ȕ��4���f�۳�p�pε��M�����E�|m���f�LHt��2��_�
y7�a��(�k��y7XB��i �q6�(C1���6��2�����zpY���lg�����s-u�����H��UB��t~
uu��Q�	/�T'�5��`@հC�a��6`[c��A�A�%"͛1�
jG�� �qL�,�P�WΓ݇3Y����/ѯQ;y��8��\,��O�N�#Y�-]Q��V������u1]������N��dfJ��0���� M��򢒳#,}�D�i�W��������ɘ�� �7��*�
��{3�m�JE$�g�g����U�˕z�K<�;��/FM�Eg�P�qW�g.�<wO��E62_uU�;mp�}i�}PfM2x�gSs� ��X�9�b�� +j�ո��0���=BQ�``&e�vg�ʭ1�i���d2D����;�~T�ڼ�b����Ju̗�J:"ui�p�	R���9�����0p�-�95:���%d����W*�[?�	�y�g���K�U��|j��dx/�Rm�	���".�����b��&�R!���tFQ���n��%�z	��҇#��p���k�CW<ip�=3kl� �����Òco�e��h�r5n�e���R�#���_�ʚ�$R��?g��U�O �1)��m0�f}I���?����k���xk6�Ȉ��B��Lck����&�Bʝ�sюt�wa�E�%��(��b���>�\9bC݇�"1�5��c�r� ����d���B�Q��Z��k\����)��<�h�&U�N%A���hq2�c1�Z��L�62NmÙ΅{��W�Hn.���_)`� �^
�{�e�8�"9�C�8
KB�����(��,�di}��W�͠��i��B�t$h�y��<}�=����GaQ�kɣ�n�kR�d�&dA�J;���@W�h �n&0�DI��c�Nbb����������C"bx�ԪZC����j�;�#>��H�Y�R�e�C���
v�4F��e-�������x��x�d���P|��a�[�x�;̙G=��>>��'sp�F�f�i�i� �R�0�H�ܯx��Qk]�F���zSzRe#�f��X��u��YA��TxZ�[7���6h(��>�V�C1��n��밒�gZ"��})^�Ǒ���ͯ>�
M�b��'���X���e��)�&,�=���l��5.1v��������R��i>���J���K��m���Ik"�ҭ����mFg�{~�I������R�J���F�Y2����VM邋h�>?.�ԁ�Fy�����| ���g��}��;e6��	��Ǻk.�ŋ@4�!2�|���W�I#�P�ힷ�],�iu��_(1h�.߲yJC�K��D�T��qh�^P�`����f�n�hw��U�~�H�o�%v��,�"dst\�?9�%RU3��I��d��$g����׆��k��"���۴��D�ց�K�@�(����Dxw�3��(w�na :����y�{Wj�������v��fR�w����+1 e����=@1�oQ��$�1U���U����Q��4��q8���0xY��t�k�D��*�Ґo,q?YI�D���j��˸qR~��2����Ct��m͛{Q"R&g�����F����MQ�6�Y�W����F���I�(sU��aϰa�i��'pr�Up�� �����s3ن]��~e���g#�t?tR~���"uP��o-�ʗ��w��h��o�]�ɌZu\	X��;�P�;�
1��18cv��M�(k�HS��VI�I�:��)ႅsO�8��7�Ór���ό7&ͣ��Q��VX��dU��|�<N[���a�]%E���F9��+i����U�Đa�i��y\�{�8��I����/ԝ~�	*)2����d8�K`��:5�Q�ݽ41�"�eQ�|DǕ�=�Jo�-���egl34�� J?~�6���F*�x����7~����kM�4E �=6<�r�I����SKԭq�Z�*�lCA���hD���wu��t�yT��A���֊��ߪHU�~m��u _Z�0��:59{�B~� ��zZ��bGj�D���3zڗ/ZRDU	��c��[�8�(!�U}H8��X$UF@����`���٣��. �  ���'Mb�,��R��M���ˏ�$\��]��M$~� 1H0r� g��ʊ���z5��鰚|థƷ������r���������C�L��`�&�]��:j�B��y���j��K۶����28��u2�{�������=�\?y���DK�{u��H�=�/��Y<�QU�5E^�:iHX����Ds���H�A�M��o�B�1�l��r����s�����ŕ�:o$����W(aec�T㑓�]Ч��a����Ծî4��������"�r�=?�mR� �Ӆ>��{8��8�%�tt���ok��؅Tw�����c>��t+�^�`�@�����B��5����fy��x���m�J�Z���3����x��#Y��W1����ߡ�mK9RO���N�ȝ�ׇ��6���*5��C*a˛���+فK��˹��J)X�l>�hMƙ�gH#�qc��Y/�Mv�9bI�������z��vk`���4���<�~ӝ�;�����p4Б3Ǜ�8�2��KAjp��z{�<|�41�+�]��<O�=_����V���-ҢP��|�sQU�յ�s�7ؼ�����4*�E8$��kIuh�V]�g3���y�%v�rS��cI�D��W~����ʧ�R�D���x��Cl��ķ.>S���N��IU48�X�8��7�CGdM��������U�t��"T-�u�2���"k�b$�0�b����C�m1����rue.�C?(�V�[; �(T��G%���}{K�.\�:��C[�W(�Y�����xѱ����)Ģ���[�������4�`O���I�Zwd��?6m����9�T.�T�}�-�kI��ܬ���J�"�nQ�ᙯ���S�%�VH��\��X�=p?v�����?�U.ژ�Z���$#e�(�g?��� �&dTo�9[����`�x���Z��a��˩�Bm���VO�ʚ�
!{��Q��Ҙ)�r��;��)'�6�S=�>zt��ݴ�m��C���"��G\0�s�=��!獔�p�"�~"_���]���%{*T��* ^t:4JQ���ȝf�=p��xo< " �^�v��ʽY��DZ�W�0�5\d+�F��`K�S����}��y@�M2��r'k V�c:L)�����gg�/������m�����S���&�k��c������w��Qg9��Ӕ�o�|
����Й"SkN�&j�e�t�dÝ�S���r
��aK�dP0)�k�}�.��5y���d\����i:��k����Ԉ�\iG=o��s�> �q�W�R;�/q���Fw�2��|`�A[��'Z,�g�ȇfFc�^#L�9�th�����2�CM�p�	c��98�a?�f�D<���{�
�jk71��ŌU�U�����B�ȁ�;'��lxT[
sE�ʼ�������MӮb��e�
(d���WnN��qo33��BĴi��O���΂{B�.?���T��_�~|�sĤԠ�N���X6C����磝h���{����M=*!@æ�%�Va�~縮`�C�~"�����b�Ab����Xn� O�����^���\��<��Q=w���z�W���x���
�:V�4�U��V2_0���J-�~$-z�N��O@��.�3��1�Q��]^����=~-RaTn�R
�c��)T݋l��IA�r[�ܞA�ᅫ	��]s�W卵!�H4�~\T��D,rW��Ѓɾ���i�ð�K}�ܤ�"��lcߣeEL��T���1,Y"D{��c�P�%;(]�+˭��[RV���
,�BYվ�\��z�9l��1�=N9&w� ��Y��s�/��s��	mn����5�yS��}k6B&W�m�TE~����<Ů�`���\˕��w�)z�<ӏv���8�����,3�
CGY��,6�:�/f����4��S�(�^<;�<����<�?�n���x�kuQYPS 	.n�18�ثԟ���gB������֋O{��/�Yz|1�_���2������8����!���V���MP��m-ld�^����dGU�0�&���/�6���aA�����~ÅY��8���={�N�A��S����]����������#	ƞ&6&�̅w��ܻ"��["ּT���?�}2|O�.��@� �ֳ�t�~'��@%"�����;qt<98��N5b)���~�����?ɤodI�Dٽ��#����-vԽ�����	U^��ړ��2�ā��'趂w7}+_�xZ�p�7U�!����/d���f!")�h0d�E��*���9�����\y d`���<6�� ��Ho\s�`b ><�M�@I�I>b�T�E��&����)^-z�͒�H�I�.lN�=��eT���٨�<�GgE��Z��4�-��nn�v�!�G+��H?k�����n�>ݹJ�Iч�._$Q�4r����m� {���e�:'����J��c�������5���'T� �9ev�Y���AN����GgꯡE���77�	:-NB��� ��w�I&�	H����XQ�дk�"s]s%�[
��H������O����;G^���u�h^o1�J�|�n|A�L�1�G~���Av�]
���I�|�;���\&he^vk���<����·Yf�3�ce��x��z�X���� _�k��QX��<�����y�3d��edU^�^��e&w�l��I�\�|�ʐ�+g�01^���B��l��l���R��4XSDQ;��3O� ���LQ�jit�����2��,�ӱL*���&��D6�����7 �0�V;����^<���`��/dND'������[���r��Uϲӱ%�M�U���	x���㺦��?	�bc�:�4&먴��t���,dH���y��p�-0췅a��ܜ<�۴.	�͎�V�k�h�,(����%�*�\3��o����Y=��������`�AM�5�!X�쨙�FO�����
;M��L�"����5)i�Obx��F{�Z�s�����7M����)"\��,�F|���߆6��ln0��m��e���ɆO�Ơg�J�}�q��!���G2u��mHEb�玐o�4��=��[�_�"ㅄ�Js�$�g�4t�G(���ACe�4k�f0�U�GT>/ڊ���V:k|4]��B�Hhrj���$'� G�9/�,�X�b�������m6��ֵK��6d<����9g�[��J��6�~?���q����t�N
�Q���ed�F@oğ�BȻ^nE���� 
@v������w�==�]��5�i��Q�B*�/�����$`�h����Y��Z�8�����<}R�à�����q(�8y����ک���=�+d�1�XS�s�Ĩ���ᩦ��䴃��t7S����D@F��ؙ�T��3���سyh�<%�$��ϼ��?�y�EQK�w�~��V��+@�	Xv���Y4�����0 v���]��J���o$C�U���7�]�8��-���H�����dWq�=˙��d�����4���X���C���}��*������n�h�X<�s�x\�V��2�`�-�kM0b�@p��i�ng��
�?����p�4 y����sWu����֝1&"��)�_����V>�S���k�x�^
01�Ol��册�L@g��x+\�c��D���㵚d�N�|�	��⫿��x��6�C���Ҭ�m=�)�;���4Z�ėdM�u@��2:,a��Ѹ(n6�J�2���Aɒ��*.t�e䦹P$x���C39D ���n6������o&
�>�(��P(��D1��mꯝ�>�B�|�/*oE�`"Y�B6��M+�Bp�®�!ӏa���[�/P�L��"�����C:��8$]����r��Y��ƚg�Ӓ�NV�U*3AߐNh�t�®$���ޮ�@B�|����P�+�d�o���������C�~�[�����n?�7et�G�tx������
���l�6�nD�t�2��wJC�̾��p�K�*�b��TT�~�<L�zIjuh�H9Wbl\p>+'��S���jiCA���p�8��ջF�g����i����cN+����]�x�䢎~�����u��e/�S��cF��c%��o��k�ӊ�<�I�q��W�,_Ga�3^x�2���.(���*I�@g�7˴xc�{���_�������OCF�Pu$��ד�����K~��[+N&W�me$B��%���0�/eD�7{�Ғ��zߑ�b}{{����ԅ�z�~��:��<����+U�٠TWf.�_�t����¸2��s��a��J���R	�ژG�_	
s�I�h�C����,�d�\���(
b�� A	ɲ�1� $�fh=_$;�����I�CP�*ݭJ�Li��MVG�#m,�,l�9�G%�UBm��=��Ԋ�[D1�2�΅��J}�/�F�7�g�x��~�I��<��Jr@ͺ��Hd�8�{m|���?d��d;�e,���5wr�9�p/4fs���
߸W`�S���7�4(�qoq�)���Y�7&�|W����1^DR����g���Z���ŧ�r~�<3��J����(�d}�"xK���J�Ly���~������3Y���),��830�
���w�
ߏ<d��+���)\��̛D��|9�$	�\;�u�Y�۹�(j���EWP�v�[Hz�s����ҁ�SO}̒Z0���*�H��w�HEV+&�U���Z��H�.}���uG斜_��BC]�m@��+C��-��&t�+����4T�3��*�{��s� �gs������s���K`������䠯�l3��P�KsD[0HQ��5𗜘��F.�!��ʿ��S��-�0�9����Ao5n�m4�����K/$O�YE�F�>C]`�6����!M�������P�Va:�g2E���r�^l�]'�����/|�"�<-�A��\$�	�:��&�_C��}5�s��F�5��K"�%u����Wg��f�ySm�=̈́���Ӗ9C�/�h���]d��U��;V�3����9���Yd[���� ����
r�x⚨!��>C)g�O�XY�!�rou"~�+�4�|�+��ufM����d�$^����E2�i��@����[#�D_��υ�5���G�E�X�{�P����e��
j�
f�#2��W���>���R������z��e�<q40��V�T�8�[�	%�`0��G���E��Ƚڎ����>�@mA�N���W��c=4b�>�9х�I/�����μ�^0�e��ŋ���0w���H��7����Ex�guY�I%3_�)30�&�Љ�^��i��v�S�Л��) ���J���Ul��[ ��p�_\���������Ў�;�ZhVn��oEn�R���@�f�W j����eG~%mnM�4��|�)�#���d��6���ߊ���ߗ��<+Z< ���M����zS|s�p[\��wL�F#�eP/���h}�������.��YW�T��]Q���\�P��\��<�d�'��ZX[�,��}+D$S����נ��B���x�	���>$%�����Ð)��G�&�5����
���׻�s?3L:$'%E��Vɝ[���]�v����J`Θ
�9Ѓ�� <Y�jqՀ�jAY�zXnqu�{cU��'zI�13$�b�S$��Da#��61�	p_�<�_�.�_\�i>y\Hp���O2�}�w<�֕�O�Q.���,B#�OפM����u�+�BV�Es�M�Zu��gK��᭪B���0E�t�:1o*	Dٵ|���=S~���Ө�����\_�k<m��tp��cT�g:�%p㛖O5�Lb𽎬��ީ�E{��fd��|�.�x�K��J����S�Vʸ��R�e8,2��l,�'�u�|%A�:	:WTh�CL�M��P|q���ۋY�Z��!X_���=��DH�Cg2�� %�>K���R�b��d�[��E,�L}��~k��z��(�ɅR�3�����7����0n2���Qh��<.U��t��)&!z��P�$:Cw���6c.��D���Ҝ�?qw��g��?��!�ğ�Շ��G����ק���R�ۜ��4�n�f�Wn���N�z�fI'�9�7e( ��s3��(�UN�ؕ^[�$�gt�Mz5{%����77�	9+�J����$��L�r�fT�����*�z[��XlxV64EB    fa00    2bd0ض���W�(X���N���o���S�&�)��Ӝm��/m�8��M����e�<��Ӎ�%EA[Z�N��#���� ��h�j�ޕ&;H�ap&
<�di��JН	C+P�<>�ЈC�\��mW|Gd@�j�Tw\��C8�Q�v/�p~e#TeVnS�2_��Ѯ��~�3�{$��\����Pu50�4��`&�b�!JKc`M4��ǃ7G
A3�,�ec}�A�����'v�i.l��t-B��+�aІI�7�/�ᨥS���(�8Bb05]�����K(E�>�����I��ENZve+a�jvl+,���(�4�%��� V��k�34Y�^�ۭS�]?��.���][!7T)�A�ٹbb�����z�aG�~a��h��d��D��šv��ʱ۫[#)�)3�@��	Ou��	/�t�ĉ`���*��SqUT9#�݈LksU jY�0`����g��+� S�����T�}��DB'��a�&�))h�6�j3�^}z�Y��Q��qQ/�p�� �x������YVG'���Q�l��:,t%gSaDa_N�N@N���UU���W.�հ=͋ju�u¨'e�϶��F�!�*6B]�};��ƢX������l!����iZ&�Y��c�3�������b������X�j�"zO2�2��=�:�5�yT=�����N���E.�<��9���?�;�FM;���LS,�KS�J�7t@�T\�gh���$Ҳ����`c:���]�FhLi��g�اW��<[�a�M{����ˇ�cl�Y�vl��`޳<~�k��J��&H�3��.d���" �{ԃ7�z&��ޤ��z�v�5+\f�WY��j�2�j�.��>J�|c�S��p��*��\ǉ7���q�I��O�?8���G""��f�gڣ�ą�FH��<.�2��şR�'��u�¥U��т t`�T���G3]�FJ�����W/��}�CC�Tg[�G)��jn\�����<b��BV,
�=_�hsKe������g��I�x^��v�@vS_�D� ���v�Wmz� ������)���#q1�1_B��N���FԺF#��CmA��B̡�c�(�07����|�AϲoM��7�v��l:�TeiБ���=�W �=��X�:�;�����,��'�1l;�|ց6r8�����=EoR�_|"_����:�O�Lib��(�;���tj^�`	~�����������*��!6y��"x���"B@�x�^w[82�N(!#�,
[�/�q�e{D�6���{%3�cZ���d�=�4ܭ�����i���m���d�l����M,	:��3s���8:#]A�Yk�s%��lk@����u\����P^���ԭ�N�N �(St�p���ӑ.�����rǢjF�T�w_��u��̃��v�J�X�rZ�ӥF+�&�_?�t����¤��k��-�xE�
�<?�f���h��Rpk�0M�-��mS&������{$���mM���X�%�0�R������e��P���5�A��`U8��u�����#��;����TIQ�w�kG�9�Ŵ�u�o��<��W>EO��u��̖y�gk�A�fK�9�R@���X+xZ�6wGl�R��#��U�L�z�p�-�-�����뭱$b��>kw��h��
���Z����kÙv���K��ˤ�w�*'0S�J2�GҨW2��8�o\�����dXnJYw�bR��@Ntk`���G_W�p��|G��C�)UT���&��w�i�,/��g������	�߀�mוR�����vuxS���6�Tՙ햱��=�O�U��n���?��?U:$gǌF�Ƙ�\�@X����o�
��E�UF+Ƌ�K1�wA-��cL�S�`	��m�K���Z�ȺS-v��Y�G��!-��wi⦇"�]L��(�k~���j�\l}օ{���o�ЫM�.��"�=�\���ʉ�[8M��c��a N���1��x2>�B����P��^�<�b�m��x�ě�f��VDDR��**��$��GF�B�`'�k��w]��E�X����0DW:����@%�e�	)+(�FY��@F�g|xo'���~. @��|i���d�nNFcvnX��qmd��e�ɜ��P0�sܰ�������;�m��ӿ�g�h�4NC�`�?<�6�������(Fߘ�Ǭue-�C˵�]���>��hGVY�;a��iM�ϧ>��k�8�d�Lg�[
�*�׬�&���	���+h):��y�鶗��J���X�>�jTi︩Q��Ty
��p��Wk0>Ŝt�43�9��vV']�>�-��/2Z,��[����(����Ís�ʫrN����NhV�ӭɀ=`�!�vt���ٍ`������Ymns5�|Q�j��	g��
��w��=�$��8��8�N}s�<1�
@d��Z����P��п�:�YOW���w��ΉD3/�^�ze~��z@�}���N�O�D��nޢ��#���+�8x&z �:�5 �h���%�|<��$��w�Տe��t���e��1��,�}��w��w+��}�(A����|C���� �|� �Ё\ ʦ6�u��`�4'U4�J��8j ���{t}�ј��A���>ޱ��P�`��}���~�s�������p�7��<
���yr�g�(�+��߾O�v9@�l�m�\���?eX���+�:�|���>���<絉5Hh�x׹
����8Ņ�T����L� �1��_��fR�j�/ԓ8-�#8-`-J �f8IH�d��MUC�+=�c�k�"%x��j����y2 �����b� H8�a�C�3��Q����]��	���ׂtyS/
zq���tg
,�`�M4`���#*�M�&��Z\~Zd6�r�(@��dg �S���{e5�&fI�l����eɫ��q`���1(;����$�	 BR�{ۊOvP	��?������i�����!U��-ņJz��`Y�]d؜��W�7h��\3��g^���,�ڞ��hN�b�N/������R�b��J(/�փ>.�>���Ywd��A�ש��a���
K����$2*v�R%�h����^&����1�Ca�kS );�)H�L92���^VF�1���jE�����Q�����	��F���ۃ;�Y-� � d��9ܫa�Mr^�I�<�#{��j�41��!H�04�V����%�7a�4�7�v�vfK}[:9�jwf��%[��{	 '��xU*��t��t I�W�)=��L#��؅Fyc:,�r,�w&,DΟQ/�Ԟ���A�(��N����?��OU���V� Ŷ^»4�=I�n)_���?����$l��)��2�-�Ʀ�l��.]H�Bstl�r_6Tk"^���L������U���D��2�ᆕG�0�6�]E������.�]w��ӿ�/B���ߎ���-%�����i/�tQ���#�v���b��ӊ" ���}H箋�)���؈��7~[m���'��,��/g:.<?U�C$�Cc6e���Z6%g�<�,��iJ�o3D\[
f2��ySC�E�XG���NB
V �L����,�7��+�G�~Z��H�^�u5��^:.ԁD����G���~?�7��jy�1��*LAPr�;ə�
���灅�@,̷�\�����P!�FqA�W<�'��Z0IE�Ï�[���|�>M������h+V�,�����V0���vd	�^31i�|�`�(u�	��+,��	P�𖤤,�g�/�v� ��ge��8tP�;�	��>�S�O>b7�B�R x���5�v��H����q��C���cO�s;�Gsd���U
�����NH�i)]6����7g�Ho�U�?�����Q�)���vI*��~F٧{$k���l�Ʊ
-M[-1���g8(%��+�J94��c����2�%*E��xko�+�`�r���ظ���ā��6|RB.D����|'+�x��b u�!�C�dB{7�+��|�G�ǋ��;~�W+
��j:��`��I�SD�]]cY(E-��t�0P^�kp�G�)�����	���I��'�$q<��#����������.{��x�k����f���	�$�ڶ���>��썸_�p��ޖZ�I�'���C�������t豕!����cJ�X�2;��ѕ���rh4E�7�w~�Qkh����=���I1�ixd$^ˎb�������֭ԩܯ��{_w�Y)�{S�D��}U���;�����Q22/�6���xݿ�>O���y��O酥D���W��2��
i�X|�M�p+��Ng�]��k����.4�>����[��7��Ӛ��PA��Y�d�;�� ��h0��a9����gE#�n�D\nRG��_�����R��txs{y
�0B\��s��Dg7_k�Z�*���?6�e6�%\������
I��_zXߝ�O�};ӡ�2�A�㻥�U������jO.lT:�m4���/��A�\���F�_*T��X]C&������Z3?�
�l�~��NH����������`���b��$����Fg�s~�86O5�"� �"F��<A�.y�~1	M��8��v�m;��^���l��&��;`]������j]-��]X�H�y��2��dE x����]$@.={�X�N�����%����}��	f����fJ�J����.s�'_a�Q6�2LFV�4���vmm��̘���dVR�/f:���<5F��s�Z�\����}	���~���^����.CU��w��P���I�A d��p6�u�4�(jlX֑X�����}��'��T\�
 ��AC_���c�QWS�T���[�������w��\Tkn�vj�,��l�d�� ��H���K�@a��bSB�b�%׉��ӎ��o *Pl����Q��Iˁ��a����Rr��m�ېs]k��0�t:��Z%���b�f�S�k���m�W��ͺ�:�`�����x:N�0�"A$�����y��k!�NclɡV*=: �ȟ�|B���.�rY���i�P�\z||��u��nM����czÀݕ�zA���Y���Z��KeZIim���*;KX��n��
?b=���U�&qHd���Kh"�HڠJ4�H�mЖ(Ϙ��Ъ�XíTC� E%8���C3�U�����v�v;�����u�(T$�AD��ݡ�ׄ�A�x}8��;\�j��
$Ȭ�x�jCSex�a?8h;c@w���Za�$u�iY�@q�����-�� ��0�2 �!�?�ÿ���E��0v��m8�,�i��!�d��cl�ö�dߺ#*YP�h�|@�,���(�r�A���.�M�L��?+ʫ�'��6�G���p� M8�3�Ze��p��7w�΢��8?f2z&�o�A �(��e�V�$a�ZJ����!�2��ԚоuI�M\�.���Z�7������M���	��z1�Uo���VR�p�4ͻ!(�H|#�6�uw�yۑ��ɩ4���0R�RFJ*Ƈ��3�H�"������"|ގ��ě�I����k�cX�
��H(d�1�U������x��_�JP�w~�\q>��r�^A�]���y�آ���DQл�M�3�Mh���i9:�(���N7B��Ւc�^nkQ�=�������"��Yco!�q�Vo|F��?�Rz3ȗ�tb�,d;ٝ�Gh, �
��BW
+�����'բ4��J��p���b1�������`yC��S֣��?pB6_=�, V�A��h@a��:e8�#�"���=���{�VӰ�ѓ���zy>�e�t��� 6�9�6�ض&��a?��׍���x��LFNƽ�4�v���=����;�<L�z̑U���[�y����+��l)ęL�цr�@�ߟv1��B��ހs��
e51.ً�`�r�s�w;g4LZ�+߿<�_x�0�r�����Y����n{#5[xU����[��ۄ ��������sk�����$��=�����y������YXe��4�wM,O�����eJ�}����ʅ�5O�p�û	E� �T����b���h�2�����᯻�� ���p�Ц��M���O�W��$ �0�a��=C(I�qE��nT�zR6�jL��:(S��P�1�҄5�.@Cv�*+ZXMڋ���!��%*:8�pT��'ǠO,$�sf���\ڿ�r�P	��R�6�3��Ȋ�Z� Yln����V�q��&�2I��_����*����Ʀ�Ᏽ��-����b"�C�=�-�˛|.�M���c�om0;�-�$�z,$�������\�9���ў��/���nx�o��y���w��ӋJ �&�C~��u���V��;�!s2�3��w�Tc�ݽ�uÌB��{tN�B��B!]��J�\����K,��;�d>���W������q�?���`R��k���E��t�����
�0~u:/ i�ʷic��o�{�E_��N�U '�|ԏH�h�vj�3TR����/|�z���tW��^��W�,?`G��!�����
��]/��J׺�G�(�w�)@s`�Ѝ�t�6�^������5�����6���k�[5��Jbii-J|� o�6W"���{�C3�}:U�3��PQ�i:���Ґ{O��x�U
��84�X&�-CV�k���
xz��V�[�KPtY���^��d;�ͫJ�XL~V�3�ylĕ���i8���6U�CbV���rw���z�����	hHy�9ZX�{��4g���u	=�>y����e��L��|e���m��ڟ@�	�~���8�9��}ث�G����}�'m�%�;u�O�"�6�#s���=�Feߓ��2�J/g��'�2��	�}�����	\R��-D��J0G��"�;G7�\�/O��� �n�`�9Gi��qy�9�a�u�j��$'�b\#�Kk�Sk��d��}	9[�Z��X��%��:�L�Y�@A?���[ʡ��6@+v50&Z��P=�Һ���j)���F�"�g����6���<�T\G��Gt��n;��I��}lx�*g���~g�����V(���\J�Y�Ln��9d��qځ��=��a�'U�L-�0Ơ]�*!�(#%-G>�؇����T.�@�<�utX\����[=6��p�H�A����8�>�Cjs�(���~�/�¦%��]Z\�6G��MI�Cw��H�@���ss�'q���`t��~jb�j��{�7�S� k 6�Ԟ;G'�8I�5���Ub���5�������g��5��9\�5��(@N���/׾��"�-��:��.j��~1FH�����y�����2TD�vW��(�K6�r|)�� ��������[�0�DX5<�e��o*-�*'3�`X�ˁ'Dͩ�Z��y�xw�3��8�e��6y9�?,=C覉g:��������e.��s��LJ��`�Gy�V��>N��"�n
�b�dP`?2\V=�oIq����b"�J`�"*�9+Q9R`�.�΂u�`��wZ��t�*�:\���ީ��4Q6��k!��f�焦���"�5AN��W�W�����n]JRk/�t-eM�o�;u�h��K�L�AY�)���q�̷eUM���Ԩ
�c����fŗoz�\eO���y��+���b�����Bz��9.�9��S\{T��$ېUɗ��{U��z�L��ր1�C(i�y�Q��J�2���Byq�3����6����\Q�1���i.�=�Gk�oX��-�Nc��T.� ����57(�:3cb_��iA�ix��o�h�XDe�Z�W7�����skc�ity�(�b����Qʑ�W�x�I��l3�r���D�e8E�\?r�t�ڌ{�?.z*�w`����:P-W?9�}����*�<�f�ߘ�uX}Q�+ m?�8u�%ʌ6�/�9��)N\�C8�UQ֒�x��w���@+<����
G���omd�ij���EX���ɛ�^�P��+'�_�g�"B��09���P8(3Az��'��ی�3� ��A��l%�[�	�x��4̘��Rt=���	͂�C�ߟk����ɔǑ���r��!��ɔQ*6!z`.6��^
� �T���>5����"���L'��b�M��BG;�w:k�c��;4��H����I���E#Ǖ����� o�"�L[JIb�b���������0�+~�����/�R��u��#��cRU�H�C�#�$DzܞE삡�5_>���@��°�ݞ[�D��	��w0[�~7�Ĺ8K��%('~z � l�OMAy�/�·�[N>:�u��~TeS}��@��"� ܺ9qs�	��3	gM*ݥ�� &}=����1-�c8;�e��^q.4��3'J���RAT�]�����Z�q��Ɇ`��q��?Ť%��L��L'c�2(;��������J�򠫐Ni�}>?�rX���ѧQP�=�-����b�[t%��vQ�a{��#���>>'�z6��?���d��w����1�K�@jF�&@|wੁ��T���.ӧ�u�-� �5��Z�c������g�	-�伬��X�QK�|�s��䅹���5�JD�P]#r�尯eL��pf+�g�嵐MwB5%f��ۤ/��׻M��kr��[a2�Pj��o��ֹtH�9�7輝�wz�	$�Gi�w�d0��7}��1ߠ�����`q�_V�D4�H��a���]s7��t�.`��l���2Z��}uJ��@����n����Rq�
^	<Q���t9��߳Yf���t�&�c����z������py��=u�	s#ɨQ���O���x��W>I�0��kbX��O���9�ţQ3B�Q�PSNf\g�C�'�Kei��.�FO� �X�m�=
&�g�P[N�Mn�B�o;����F�W-�
�2����/���QqH�1����g�"߰tu��f T�.���N��:� �tjX���������]Ĝ���e1l[:�J$��V&�1ǦB�����?��'`�P�A���������yƌ�|!���E &m�ߞ,ւԅ�~��V]̬�(ebŧ��ʅ��%�/�����/�1k
1��$"w�^�٨(>��z�*�XY����f�Af _QH�Nբ(0�Q��57��m�H�A����3�E����m�(��M*(S]|�˙���w g�V�{�d� �̌�@�,�&�a݀/�hL��\�%Ŭ��[���7'�t0:�������$�b�b���FC��M�)v�DY}�A�%�|uJnΖ]��o���q2�!�Q��P�L=��^�:w� r����e/�_�rG>�uNԔ��gǊ��&̥�DFN�B$!Ji�v!�P���	}�Ct}���_��Ъ�4Ͻ�`�A�"^Z�z�E�X6�3Z0�*C��z�Ѡ����׈	%���2
y|��ߨ�!��e�|N�b�QYG�N�!����TbC�ؚl�NlQ���������^hy{6�\9D&6%KI�	���� lU��ߋ8#��9=�3cG_�]�3�P�=��hLg��R���nد�j�O�Xc�2b�2��\��w^�1t��$�L �������؊hbp�=M�gg���w۠%2rJ8����#�6�)��峡Y�y$���Iu��w�U#V�c1/�i��&g�?0}%�:��=�Rzh.s�Uk�!�J���*��!�)b*�o�1̨�?Y���d����ΓD��'��-����������ߑ�w�jxʱr,�<U�]l6�]����@�/�����G5)������ _e1�d�m[��d_��!
�ĉD���둡5������|������3��fAW���k/�����:f7���1!8�� ���p��2�����'^�3q�Z�1<�Jʜa���mr�Cr�(��K�ThKc����|&<�$tfl���3�X+�ޟ�n�	U�Y	\@���|5�9f=�vaj��@������7�0`���ʣ�!���He�7��j�Co
�r�V��Q�	C|�)����=X����I�����2ݔ��<*�]57�Y@����;����Y����ཊr��O�?#�� oɿ����]xи�m�cY�p�~�->N�s�z�n�B�4:y$d����/�$����Eղ!�6sx�$)��׊�����B�.�� 
lz��wu�_����	Ҷy[`<ڝ�**G\��we@A��#�4�e6j�<�HU�Zl��a.�8�/Y�	y�eB���k`w�[�&�Ȣᙆp�����VE]����q��ә�ͥ�ծ�	z�[��Q���.�.�z -��ˇ��t�1糳�LL�����Ւz?=s�{į��C$�M�F*>iJ���۲��v����u���n��|��[d�~8��D���t�6�"�:�ƫ�|��>�X޿ڵ�����E �Q3yX�;C\���
*gnB�is�t�z��{Z����M��r�P6�o�D}�d��ŀ_q��'J?�s,��'��e�/x�*(:���BA$��B���h2Cqi�|.i�S#������e4�ɬ�}�
�����v�^�`}]c��}&A���-.���b�`�S�V��������� ��%������'��y�O�ϕ���͜��S,�Yy�e{�j�K�@blڛ+w�F�A��Dy}�B��:% �dYv�~7S�+���T�Q}�x0��s�\	�ъ��
�]�Y���x]&۸J؀V���a�z�,Hoq1����C_�JCR��oU(�X������"3=Bo��s��a�GT|�B���Q!X�_SG���{�����S�$-��v�)I��9����n����)���/;pz���kS��U6'�����[��cYǧ&�9)�D#&���h�P��%)O��)DbY5 ���8�(��ݳ��?�ͰG@1~�Xn*�Y
A����t�8��DY`�1f[s��5
�yB�/��+��T��pڕ�C�#DM�#ŧl4��~3�ڙ��H��)�XlxV64EB    a2cc    1b60��:�|�|y�16�/�n��2�	�F1��g��r��	&������� 	][R٫�s?��Z�[p���l�<
�s����eI,���+畬#�z̴��
ۻ<}��mV�T���W�%+���	<�/o=�@�B$0w˴sC�]jH�Q6�+v	gˤ�i�V55�(y?"z�{��-�Y����D������,��,D@�I�t���P[ꭠ�z�M䳙ZS^�X�cwo� N�q���٘�>����jG�{F
���c�|���I q�6�q�������0mZ��oꂅ��O\(��Ȕ_����:�t(��V��F[B�s?8|�	"�1�Rf�����r�k��Cp� V�C�/H��s/�/#C���*X�]0�:���BD]<$��dwN)��/�[ٹE�Ջ�Z p4�vJZό����C�(4�7�e/.W�|,	�Д�����I�h@{]'ך�~������5&#�r�_���jo)��������5��-f�Z�/���a����>��߸���Ҕd���C�ɝ�J0���G�~r0X�=�zYZ�wV�l"�/O$��[s�O�ɜU�P��1�o$����E���{NH��"�˙�ۗ_���/�f��o���,ӷ&����(�X)V=6y�+#�E�SyHM*�����]S�r���N�R}�_�B�u����������|�ct�K#��S_8N|#z��E.`ʛ��2u�B�6Ww-�pkXt�m	y�=5}~���-O��nH%����&�B�-1�#A>�TG��Γd��ka9�tsE�~�֊�E*�!� �����ȥ6�����MJ
dd����M��w�
YO�1��h�5Bv��+SS��k�~���I�>�.��4�Ԧ�<�`��6H�p����\F�|^!�����t�Lq��@@jx[0Lt��L�P��-=�0�EȈ/�ɨ��vΨ��RH�X�.��5�����7	�+��n ����R��7>����\�w�Q�g-[�����?ufb��ڰ�4؝�xj%����OnE���pr��ok���r.��К���gWL���^�B����+kT��bS/�LG@j�\��af�Y�����e�9�I��|c��m��t�=��?hc��X�j�7��K�W���1	��!���!�b#��۰}4���t����y�-��q*`���虮	���	��H�E�JP�?C�3g�O��DIu��r��.���U1���c����W�2��yNw�A�OZh�F0�Y��|3�-�A��h��"�K���؇ +KZ5�W��w���L�i�gN,�^c���z�+�{�ɠ{��U���ڰ�6��ZM9�]���J�x���m�.�8C|���[�E�4�!�h��%��/&�UY)��L..l����uyS�F��q7w!ʝ��<9`k���!���}9%�M�8)��W�Ș��
���~�hSU����M(D��D��y��s�v�K)��$������A?����u�3���Y�^����*���(�r&S�>��_�U���䄋1q"���Vi�u=���AH���*�(�r�|o��B�������[��skӬ�0�B^�����"�757���(��^P��n�F:4AM᠂�s�"W�=7�G�+4T����59M�ܾ������LW�������Wp�GwW���l���3d�Q�z@�����°������4J;h��}��6��"�B��+}k�v��� Xb�)9ݜ�I�������> #zl��~%an����9���4z��M3�R�����H��?>�9�w��EI�B��c����Y��a	�	��#��/���w���W}���T���!M_x�`'��������s*�K��j�?�r��<�@��|:�p�1wE�h���$ ��q!칓�d���1ʀ�ƎH-�ɒa��NC�<�Qv��H�i�Q��'���S��ѸA���g ���W��呎c��t䎧"��8���u�1��2ˍ�~�J=Mk��Ơ��`����\z��B\|˸v���C��~{��85��4�?/�VuO�g�I����ܥ�q��M��$�p-u�<�+�e��X���xs!+��&��$~�Xp�������S��;UL��gJӹ���/�x�$8ѼPo�|Y�9�*���e>�U�=1Ygϕ���m6�!2���q���P��*�Q����Lv�
�;�PUf��fn~ǰ�����|����&�[a�5�2_����swT�f=�Y�C|�0ŚB/P��$2z�'�M`6^�Y�b����Q��u�8 ��� ��R@�hه�Hm]����)Z����"8!���^�S��$<��AK����g��r�:��. ,Z@�Ul)Z&n� ����S���"(�~=Ӥo�4ukŧ�H����mO?��B�%YB�D��lFrUSC��s��P��{�-�-���O-��A_���-2�z^b�n��Iݴ�ȓp����َ�%�|�%�<#%�]��2����ŤV�����x��ғ7TZ�{03������M� ���̳���1��u	.���/��I�GWB�c~X��Y�����UE����v�s�
�_jㅋb����Hw�����&����ܻQ���BI�2�v�+a�$��а�q�@�͈?+���|Tp7�����WӞ沌����Z����sl'9	��͠�.C��a��Q)��
�0x�T���$��
f�=?�Y����uq���;�RL{��Ÿ��?(f�D�{����hkW����a�6��~�?�T��xX�<L;�E)`�$����Jzi�\�k��:�­/O�२j�ꍤ+���X�B[����z]���[v����K�(������25	��P����|{D���Ϥ����}[D�^��$gRE.�}H�e���(PtO:s6G��K��4ň�N1*�=}#��Z%}����)���32�^L�mM ���ז���#�t���l���"����[�
�s�r?���B~X��5�J$�������b�Mމ_�a�|�_o.�\g�+-	)�l+-����~-2z�����xKE�讘��� �G8�\�*[����bmG,B�;�a�ʁ�4��v��b�� ��UG�S!��%�����y$�1音�y�2��/�Q�}�`]11�Б�DsX�k=.�<FDwqքzI��T�%Ɩ;��	9g�O�#�,ԡ3��[���,>诲�j�����W��Q�br�9D�({>�6
��(j �"Ȁx>؃���&�pa��q��u�b�~Ӹ�q�J� ��[�؜&	�=nmq�}�fDK[���ḧ�:�D+��n��e�Վm{IB:�?�I�\��α�-����ń1.��<�F0f���=N���#��.*�c�������W��N�/(�fr><`���lZ��N�b�A��=8tj�:�R���R:�s�a������Α<g�nŎ.��⛊�-X��/��d�����[���F�I���{�nH�RS�́�N� ǅ�|<[��E_2oeBn�`I���Af�5:�1^�
�O�j�O������¾�̞�}oT sk	,���吧�D�\u.����Wa}89E�:2,G�F&FV�B$ˡ�l�G$����: ;`%��yѽ��T�t�,�ջ���k�Sf����B�����0�%����K��-�C$�(�s�$���N��r#�Ȟ檮�hX�/��m����FM�wj����'=q����`�+=� H�xDCCwڢ�%��'ԯ�pRu�s8>_��r�"��[,�k��t���X�^�i�,J�w9ҍ��A��y�y���K_�f
��ߏ��P� ��?�b��of��#^Ҟz�r���G��q�����k|�@ε?�v�Ez�`��r��sZ�]�W�Xx������٭1���C���h�������c����B��k]Jĉ��9ƒ���<�)�	-�[]�'B���H��qC��m��"Z�6���eJ����D-�?Y���VN:����3f�?c�ŧ���U<�w�H��-<��C������K`���TeQ?�<PD���M���X�6d=ה9�q5ډ��Ia�S	�.`���T��p߼��h�GF�7��-/�f�¬r��VJ[�ܧ1�b)t����{-I?��9�9vn����&�Gr������n�!<%����8蝎;��h�ьqwV��2�xk�����[�����d�HI�mD����YvY�����e�vpA�L���+�FT��*��%����(�R��%��H rHN����5Ү/S&E�l3�4x��s�#s ��Q�]u4��vg�ii��mՕ�־�
�I��l�'ǝl|��z���2"]���gf�8m�%�M-�+RGø�P�\�TȜ��7r��Ջ�2�Kw�u�21�D���$H^!`{P�4b����( D�5{PY5���|�I��S���N����iømˌX�[���%���x�ݞƮ����0M���@�	��vCd�r�/��vU�h<)�$�r��sn�$PE����X�G%ڴ�I	���oa^*�4du��f_��Q���M��@�����'�c�<����HJ� �@`k��:��6N���
����'K���W33Yؗ��`Nt�!�6�ǌ)V4�*��C4v��5�	q�ߑ �9��Q�S�!`�Q��p�J�|���!F��C��g�1�Li��E�������\sn+�mzZ�s�4�����<=�y�lG;�+��o�!դ,wڞ�pP�_�;��j�˳��0K� Y.@��4�S��Y4q]u��8�­�Z%��U�u��������4����2������>��&`!w�$f��"�4\�:��Y�c|��Q�N`uy��5��}�~�X���s���1������̈)MF���`	!j^�S+�A/�l �T��m��iNe��{�Cs@^�2��B�G�Qѫ1����=�#k�꟩�����5>P�Qv�N��Ƣ��1_Ʊ��H+ćK���'#|�h����}Z�P$Z��E��8�1�&E�{�ͅ���Td]�������#��f���|ǿ���@"��d
�y���f��^x��U�����ˎBɺ��X'�N�=�5{�w'YX� fi�z��Nq�U'b�:w��h��߲��[�T�m����Wn|�"jCͯqm"��}�痰A:��ԧ��d�j9F���՘�+���}�(7���/+
�|�v��^�V�L#�f42���>�x�Mu&l�����h�\nÐ�uk���l($��hKJ0�����c��I���i��U؊��A��d�1J�+'S�+�V#���xX������lJ��7U�QM�b��Nz�]�pD�>G��jG�9���~��6_��5�/�������ل1�,i�/��'�XC��Pw�e��k�6�竛�#MZM|=Ȕk�]���Bm/�pJ�4,����,T	��v�1�]w�Q_�B�:����6L|��x]�3/:�W��ܙ������-�֑;aZe,;�&n��tϴ%�A���l}�
��[]��<w��u銭�ʰ9�m�p�/C.�\|�Ù�ػ}JX� �G.Nۤ��yewr��t���z���D�唭����}�`56���6�]�Q�UA��Nby���Fl �D��9Z^+BRL�|Z������K���u*�k���~��0�h����~��=H 8+�x
m�>����_	z��TI�3Ή�)8���&Q*�G�}Γi[��t?�Qn\�?+�Q	_�eU�ާ6��~=ڜ�Z���P���@$.���vA��`\����}���.fż���V�GM-��&����v������U��P2,�Z,cA���+q|��m�n��4�� �*��PA��5sdƯ��6�,�DN�h�7�_��<ik_�1�g�8��Y��,سi���MW g���;~�N�a<3�S�1��
3��wO��|Ck�������MC�ކ����t<JqQ�É^�Ц�X�_�bؙ���L.M���/�X��o���L�$�J�)5�>� b3!l��L��N��T��0���1ݼz��b�O�H5��%�	i</_EP�+�Mi��\�j6��!\��)9�5s���p�j�����I�RCµ	�!��0��iЧ�tjmݲf�X�X�zi�T` �.�J��>ap��QL��,�W���f{�MQ���-=�޶��/��'|W��vj"X�E�\���i͓����k����R��
XBo���[��B7��4���x��7zP� $
߄���e�	�T[��¾n˅�t~�(��[u�܂�Vڐk�u������2�;��)�{�$<}=�1!Q\J� ��|թkf�.i�%`���k�^���<g�s��F��m{=��W��}�4�`+�)β*W�c��㒣S@�w�4��U�WTHm�ߗ�;G��
�Z�h��/F�xa>/ʳ��4��q�����F�B�ͥ�{K����� C�NJ�|6��E&Դ�j�X��9�yn�M1'���8���
>���U�Qa�~��W���ޔ���)�3����+��ٙ!�F�j�gi �B���9���j�^+���wm�Z�e4@�cC_��x�wB3�����Xgq����E�ͯ	�Y�A��5��-��(��������9�N��-&�J8���m�[�(<�_�D����=R�������U�ȴ	g�k��qoe�ܬ���Z��|��Хg�J��q
�=�Py�fr֠�NrD��B|�),�yD��L��e�,��k��5��cb�rC��ī]�����m�$����w8n3rt�m���O���M�u1����/��