XlxV64EB    1e92     a90�@}�ܡF�O�o3L��r;�TMӠ"D�#�o�E9 3X��md�/�&p�k�z�S;`�?k_('ܨ���ҡ-0�t�l���-;h	��J���6ױ5�~/1�)���=_�PRL�=G�YN�NBNS` j�{�����)�B���ʓ��H�H#�A��R,�4eU�50�$��
+{��t�
?�q�wT�b�g�<M��F���b�Ҟ�%h��-e�4�qZ�^fC�hd`�&�t�s�9y�jQ8k�N�P��� fj�$z*�6�}� (��Ok�#�gN��%zM�7�	e�I�G`��nJ��Y�w/��ZJ�)�y�&�$\yB;OvV V,H�Q��A�W=��e�t��{R��HMQ#���8`�u��A�ߺ%Cu��v̴���K?�^Ɋ��ޫH"akJ�lC&�����)5�[������s����LE�0n܌]3I�l���T�(������U�R���}�@�)	�"W�o�~���A���~0��i�_F�o!�b���k��^�ݓ]�9B�`�\*�i�a�7,T�D�A�3��c�Z��eW�0�Z�B���;��� |t
���G�*�B9�,��������%ݦ��mYtCX�t��
2��[5��#���Kfr`�t̂���Aj���t����2Hffk5�#'\f��xM���m$�TA��x!�%������Y pY�=j*�^�a�T��E�D���,�O���f�Ze��Y�S��B�.+F�Ў ��������9VShbh�GH^��@�4�E"|�,����ۭ�=�9��F��U�+�R��"�
�pZ�� ��
�W����,���z�j�)8BN��V�YU��5��P��&F��d��+F���k�e��?����K&^cY:�Q%}=ɂĽ���Vv�-�e`Cu�� b��Y%*�]�|���T���h��8T)ChI��\�����b%�7�57`\$Z���^�g5/�/ʹ{R���[@,\q�W[��{��!V��ҟ>?�G��;��7���"i��	�Y�|���sV~���`�b���5v���X@�a<�r7�]a��C�v 6g��n��T��O�'5N��bbf�
Dl��H������&����o=��h�L;G�!S�U5S�;4�V�e���Yѥ�P�a��n�qJ����ܻ����H��=��{�^��Ȋ��q����D�������,C�EFZ�m�tPZ�-���i|&�O!�=z"�!I=��[{=l��6:�z0��4Ҷ��Ehڤ�5�)F��/
�w��e���#F�m5p���OR߶Cw4Px;�(��I�=����C����Ĝ�X�P����2���I�c5\OpM��d�J!8I��Y4 ��7�!���鹦,�%�B���B�Ո�D��G_gdE���ޝ��-��/�����UE
�;9_)��I<�T��-E0��Eۤ�!����;�=�M��ݟν�}�H��N�C��Ft�I�ˣ� Vmp_#|2��� ��m�{ &����1:˴�`�i�cs�dASg����Y)~�9�`˧�F�3̌OL��P��5:�%�9�I ��������br��C&7h��b*��H�v+U�@�!��c�c�K�|#����c�0����^?�&^8���c��r#q{�����1���.�9����z{�P�"-M���u��>eOk�An�2��Ĥ%U����g4��4�[�\.��s�V	tS�TLw�N�Y
�����e�
�PU��I+��@�e�d-��P�b�[p�*�=j]ȑ��@ŀm��6�NI�s[S�����	��@*�����߿oa��rm-Vc`���_�_M@*V���9��
� �!�c����hbx��v=I0��o/r6��o\BB�����0�w��"(��L�?-�Sn�s�F�q>��|̼v6n�H�)��[ tk[�W��r|��aċ��'�<����E�F<���T9�{��)A]��z��}}�-Q�+��bi�W��ۈ�_{C��5�(�+�q��TT#������Ʋ"�>�sEE�ސ4BL�Ǧ?��f&�a[����)J��䤍�_��aӠ*��ld��PĹ�V>�n8���Í>L�y��X���,�z^
��%�l�!��4Ƃ[����k	�.o�Hp�5�K�R�^��31*Eł�	,A���Wm��٢�Q1�_@�~��~���(�^Z+�����D>�m��@<wY�6�&[������FuWtN�2~]֜>|��C~g�:#��`���|� ǡ>��I��$�ذ�h=!��'�q��ds�r����6ꥴ-�%U���Q�.���i��$u������:C� �w�Z+za�e�lW���F��s�m��0���n���&M:��r�[x�ju�֯9&[�E���2��%�NM�������!����)�j�
c�\ 9�Nm���?�K�¹����&���'�y��q#��%��6/�K��c�ЊkD@�G�O��\.*�M+�K�e?�n`���ٽ��fǄ�gh����]��}n5�R�yR���U\덗�I2t�;�d!L������a?�(�hrK���7.L�|7^DGw� uZ+��"���yӁ�,�� �"]���/{P���&�+r,�1b�{�v��m�`�X�Y���