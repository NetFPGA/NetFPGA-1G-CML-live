XlxV64EB    3820     fc0[�V�3�3LO.��l���%AZ�`���mmB�OOf���LX2�٢㉦�6�'�e�^#%���|�{Cn��0
��� ��:���]��ࢫ-t��������� ����LP�1�Z}��3��떷5�?!�����-{d�K*�U^�\���g��] �d7c8q*܆M^��\6=�>!T�N�v��Ot
D�;VN��`�Mjڂs��jhby��t��U8�u�_�<S�0zD�U��7/���2�O�������BF��xf`�_��W�������� �U����q�a�2�La�Iܸ(�-���g�Y(��(P��1�/!{�E��pX�7�G�7�P��*�����f����S\����W5�Hŗ۔(/dLr:񫣴����8B#�:ȡ�"\�%9ǐ��F�cvCi�j <�����i��Pe�����s�[��������"���̰���'�N{�RJܐ�g¥���ɘ�R����_�0�9_�N�����#٘(��Km))bA*嚜�!�E�34=-�!�с���k��-�ر�����8�+� �Z���#\���㵘d{?�/��׋���rq�P��.1���8�98�~�A��zI���p�cé���W��:�T��ff����S[c��x�Yr�<�s�1�k�<��E�PxJJ��r���[����ɗ0v$<�/�E�;��*TQ��Z�f"���3V��W R6.�k���ۭ׶�"&�7��m�1)��1X��4gҏȜ�9.��sZ �OX�s�����j�I�5�+?�>�Wh�7h��+c�L���2���K�h�:>�����Q�<�V2�>�q6#�F`���(փ���wxs�k͠�٣��]�l��znK�����WxE���� |q��m�6�~GD�2�,�[��;B'��X�O����f���F�J)��E�yӎ��@$�؆n[�zסr��J���þ�;�dt�͓���?��x2|v�����+ِ���H���n0ҴX�NԏcҢEr�E]�ig�΀�ѓaNr4Q�̜
H�|�c�߱�88����I�ɭDJ�e�,Qb�xؒ�FA4���ɱ��0���vdY�X����I���������o��ۛ����f~�U���;�Qܙpg��8�끧���W"��<	�!;��>����ɼ��R(��.�	�~�&_���uȤ�������ô�$㳶W���5�Ҕ��.����y�ZՈc�������{+��������M]�M
��m	��L���X�����酵NE��x%d�f�l%K>F�92�.��e|�y�:�M���q�����L��ĿTGL���b .�-FA����f)C�kPͲ����yt&0����q���	�F�?JV�3S��NWV�G��(��p�)k ��Ν23�@K:�z��{�2���,6�[�XJ����e��Xx-�s��+�C�$�J�p<ۭK�������=��<@�Dr����[��?�v�D�XFv����x.#��v:ˆ(��ε=�DYm�����|ƦY���)���?��U��>�Ij/��˒��	��Lּ I�wfʣ���'���t��k�z\�W�ԍ~��_'��w3�\ؔ��S6��1sE�Uq����0N���M�7Fx�S��Sl��rȈ�^�1O�4&7�pXI$��6By��Z��k1�E�+�DZkl�zJ�!m�q��u!/&�Bt<v��������
�S�$�w��hބ�M(��-��W��0T��,[�]7�0E���Z-ꤰ)�[�R�;��ggÓ	��8]��2�W` �,��I�l6���>T7�pzG�'?ª��i���E�z�`�F$9���K��l�|f�0? �E[�2��4߁
\6�5%K��j��Ò2[7�\��$L�D8�<�f*�=k�K�V������4G�K	��̱��vP��칚�]yu�,G.WI�T���8g/�9=0\��|/j@�q��:]�^�{�څ�����ڮ����:�d��D\���s��	k��F�^�b7�V�;Q��^+~D����� �����"-�a�E����[Y���J题����ي��$��`f�,��
70!��K���}�Q���q¨�(v[M^�K����siM�g#�ӔhR,�Kuq�ڷ��z!��=�^����B���H�2ϐ�ХH��8j_{~t�?.�"h�T�8���";)4��?�����6JxǃKۤঽ�q*H�_����𺿼�S�d�9���V�â�y�$�����ڱ���l���;kP�M�?;��18����]�nɃ��M�Û�/��=(���B
��x�(�*D0�a��"A'<�`�t)$��)d���W��ɨp���C>�i�gq)L�D���q{5�6�ur m�rѐU�K@�׶56n�4:{8����|;��V׍&{�//" ��еM��GրQ_���TV*=�!�*�wWTێ7]'�w=~M�j�����X�\�w\�/䦜�J�.�L�?!���5��.<���1�XnsN��x��TsF�t��L��Q`�=`w��,�?�ae��˫ r�����/ݘ���������⃫�L�8��7�XT;kvr�<�n���*>�i8�P�˓JL2�dϻ�X����9�锫�o1
�#R.�=($K�OI&�nO���. ��>���r	� ��0+�X���1�S�p�B�AN;�DK�(f�{�Y�}z`�PP�<�9+���|�/9����/d���Y�1��./���������)��5,F�	p#
Moy�����l�>`a�+�:(þ��1�*y�)������ ɱ A�{��spf�P�a�W+���;�kޒp!��18S�2�i����Nxᒷ��6oq��	8�m�z7���VY����ھơ�Tt�� 4�@����!Bډ�Ӷ�w�K���|�~��c���32؛���P?~�_ާ;�p(�|�CW���SW�L>6��LL���^�MO���:[�O�6�[i���fb��r"��yM�"^?��?$c��\1{�����s�s����'�^ߑ､|gS}8��aF�ʒt6 �Ȃר��4
`̍ �f�Q�.Kҳ>�̰r\��\��J�E䛿T���I��m�)C�z3�A��<����WS���*1�L�a�.(��B#xR�T�>Ő[*XY)13�&H�Pڦ8Ѡ4�l ν�.��T0BGק�E��˂r��RO�n��z�ZXhZ�J�P��A��f���5�#��旵"T��H�f�%�/bjeۼƪ������ve��X>|s/��?o���6냋;>T�����*�X8�SM� ���ԝ%���b/��4�ƛ�Z/����>�T� ���!@z�D굢s�:|87��t���z�bևD?'jqTV�Wo8�#*���;,��M��=~��@B�k�qC{����`�]���}������]ă*7l�B����� tya'I$��${�--Y�$�Ix��3#�MH2`�T��D�!5��r\�����@\���]\碙�ƞKL6�7灀IS��'���)j���6{{�)۶��lK�(�Z�R6%J���{�r�\�bZ��tg�	y���I�q�Y�m��,�L�br���[&��#]��������U7�$���<A3Op�Y�i��vB�!`U6p���}�M�V]������$(1	�pYB~� �F�4�%,���+����pL�Iq���o�X���`<��+�3%@���]��te�2�����;^e���b�p���(���������(Qsϭ�\��\��>�eQ�l�٭"`�ۤnny�h��H*9.9&��+���ԩ�]L=��~�9c,4v8��r$u,_y�������0v�h*���	5LMs��	�'��[+W�͠�,_
�\U��By۩���:�|�jU[8f魞�[��=i�
7��