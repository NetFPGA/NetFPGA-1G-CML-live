XlxV64EB    32c8     d40����vw�+}�v�$y؆��Ƹ`Ő4�=�F��)V���s�I�em+�����Yg�~5���[:�V¹u�ޜ��d�E�����?_Wj�/+\�5�����L(i�w��8���L���D�ҹ��^Z�d��李o垪k�8ǡ�(1��ﬖ��t�~M��fGeY�\d^�#�!�o#@�xQ�;-���L��!��~[�,�6!R�d�Я7�g�N���H6�a)Mi/��W�bX�N*+���� +�2�^������/_�yX$�U�4\MJa�����d0(M��w��U�}���7�K�Ίb�:n��C�`���$�	�E�Qn��`��G����GQ%�|��ԭ\TcC�ˏvЃ\h�14iV�Y��#(j\Q�����x�\a٥�i�5��u8~�鉤HeH��{������b��Y0�������V�5Iߥ�6ׯX���7D8�JK����qE�Zេ��,1���0�����Y��8�ڼ�Ia-�[�째�#����E�<���n]�5��.�z(Z��/+����z6�&,*i�.�nG^�6��yW/��@5q�S0�Mv��Fme�v�j:����VE�[��%_��� ��s&��=�pQT*/�.˗�Oq�&J����~�����{�\����^�$�#?̾���,Y�ZoVή5%�o���9���*(iu�u�����H-�a3E��B'f�":�G�|X�B��$p�z.�\��7U�+UѦ^�c%��;M�������%��Z�k@P�P�D���[g D}z�
������(C���nZ��s^�mոN�3m�3Y�(AJ��ǝ�%V@��w�K�u���|X��18�0[#X���X"��TYiH\D>�Qu�����0˜wu���m�
݋ZV0 �mGY5򉇽�c;o2����Y��S����*�td�zm�Q=����+qʻm�ܗ �6��[���V�����p�T�'��ou<��1c
a��p]��i\��)� 42�_:{[Ik#�!.?h� `{�;�����Y[-��/5v�+��4U��������@����3ƃ8������a׫�`AI��!��Κ������m�>ZL�z��X�ɘ��X@#��k��H���֚&6j�Z$������_��F�X�Bdg�Ut��;�Oc; K��x��$�P1���e�H���ӆOL��@z��9�J�`*n�[�HhYH���OS�0c�����dn���S)[�H��{�Ht�$S�i"���%���q���y�p0���pE��M�yϨ�U�n��S6h�%�ZW-A��G�R�A�*�0�����.t�.��t��_F�U�08v���n�#1L}�6}[�e�.�\�B~����N�Wҷ�d
�]]|y�Q�n�	:/��9N��	��ӧ��/R��zF��'RL'�o� �|��䶕]k,�\���o�m|��������JR��<����=M�45��#$�����<	PnRz�_��t@�Qg���KK������Wu���� ���ҥǝ`=����ƉL$��Y�Hd���Q��a=,��B�-���iq>��еz'� �X��Y��C��J���6o]�X�:h�>�N��G���L��#NՋ1͸��=`>
G�GT2Fuo�-����k�HD\Jͤ�TQ�8S>��
�98���i�^ŪM���$��t���%����k�v�х3.V_�����W��i<g��ةvj*�o�n��<dҴ@�G$5
��2����79��QS7����y -&b�b/���fa
�q=Չ�F	G
#��/Иy���3*��`�e
Ȅ^���8[��/4���k�`�AvAs�|.ޭ��W�]�>��9�$�:�knlK��oC���ό[���n�7���H�GL���p#��L�# ������Z�hVQ��_�e.5�ʪ����I`�}����a}�����ӲW�>�A����J?��mw`�bva��?0�����]6�}�>>���3�*��5�8�� f's�u��G9�z"�
 :}���"�9H(��X�&K���K�j|��8���gR?��N4�zJ6���+�-Uyܳ��KOu��;��O�U�L;�#�Χ�:`�7�Tf�o�E����u���, �Y�Q�1�9�%������c/�
�]�!ɀ�;�L�Ue�&��⎚uV�`�5�95	ff�sSi2Y��Y`ؽ� qِ��2������,���� +a�Je�r�2
rR���q-�)���x��(f,cO���Y�<
~��P�X�9PC��A�9����Fl�v_�rp��*�����^ô&R�%W�N��˥�=Z��p�-�ЭW�J`��x	~�|��]z���V������wǅ�=�����2��9=t���!C�=ύ��᪆a�?z��?���8�8?i�$�n�pI�4
�o��jR!���b�λ@y�^��aX��n�A%�b ��?pO��~Z̀6Nī��3�4UT��s{��G���FM�Z}�'��n���\��Ij/��	ÕO>�=����v�9�F�bKR�������_볞�@d�9���X�q�/`��B�`ً	 ���Vy$�I]oCiaK9c3 �[�;�n�b<8�=��G���
OQ����M\� �[&�?7�2�3�/��,���Q��#1�b�K�k!n`��x���HpD�x���+�\�li�0^'@䏝T@�����>SJ)��M� t���
zP,��ԉ���ǵԝ���(���&���.�=�x N$} �H��V��=+�����("�W�u��  !.���Sw|��.:k���D���%��y(_�4���A�J#L���]#D��Mh� �w ��,��x]�`���׳,hk6�H[\�4)Ń��J�-Fd�Q h�w �R}�YsK8���_�	��Zr̲҃�tS�^K�LAm߫Q���2��dIn��Z���ʉ�"y�q��l�.�q�XNb|�ʻ2���B�����G��f��e��(qat5�K7x�߄9�C04��F������F���٬TC�}F�@̌ȼ��\(��:ư���6�ۭj;(b_����H�G�(N&�G�z�2]tC�@
�壗B��$�&!�I����������"���0������I2���4
a�ƻ-��I7��H��p=��S�n�P��٩��ߴ i�1x4:�������+Xo3���-7)�����;A)�)L'���/��S�z�|�	�e��i��~SH���f��H
��
���