XlxV64EB    88b3    1c00�D�k��w�Ro{Ş��� +^�A+x�����ؑU����q�T����|���m��eI�C���2�_O�.͜<7���zAnRy��AH@MDl|��\{8�!�~Y�C�rMpdDd��µ�+����'���i��%`k@-��ז#�Ϭ��%>�B.�+"$H�,��ӵƔgU�>ID�'HL�O���^̡���\v�ߕ�6�s-h�� ���5NQ�����ſj��A�iSy�"����&��N�����GA��7i�o-	N��QG[a�� ��='�hyIun�ӛ!?D�ˡ��Ҩ�()��$JSg򎡨����vf�-˾'�V���εđFw`Ņ(����L��R�ȂbG�ͱ^G�-A�\�|ufc�@� ���/Ҳ����P͹ IhU��u�A�c.�T`��{P��C.,����#c�ҫu�.ֿ%���d:���S���E�^#]�G������p*}�����
Z�:x�g��^�oc�)�%��N�:>�!]�ql�I��'���Q� �d_Ӱ����t��7�V�N䡹���/�1���l��|Jq�N�2�R^��C}����V(��-�m�=��nŋi���=%�.��NvXf�ۄ\�b$!l�2pKs��� �i;�P�:�U��t\�x~��hs�Ee���Մ�W��'W�l^�a�[�+~2�G�����	(J��Ϛ�ڞ��Վ�?A��!I���ÖLf�Z�x0�Q��F��)���	�ܦ�C�ҏ�������Pa?���ݿ�_����->=�������_gY���$�Ѹ�j��_Hд/�fm�LUH>��@� �Wa���i߂{��ڰ5Iw��,reAq;�gMx+�K��\bɎ0Q�i�
h��2�@i.P<�_�����Ά��SǱ�l#��_���S���'�v�3��D�����Y��a`˾mU3}��)�MŦ+a?I�xu6��]���b�t��w�ʟ@uU x�`
���u�*�Vx���OB��)�+�W�H��5�v�hQ���TJ��Ѳ���:ir�٘�/��JA��+��!Ĥg��^c4����+�f�������B��gD��m���H!���=��xD�L6?��b\ѫ�\1�אݘ��s#�D���@�s&�����c��@�D6��D��ę��)��4%G�z�=«��ŭed{���3�J����+d�>�-��׹^�-�L�e�=����C�0�h��)!B�O��zqF"e�0!��Ok>�zQ[�g�F���N%R��z�k�
ȫ��P����XKe.�1wo	�m�a�H�e�;<OR� ���ߝ*��������+P%�4De��@�ߐ���;]�j�Gtc�))P_�:������ \$��ۍ�TY����F�>�� ���x<�����l޹�H�]s<��#�C:��"``����SP
��`5��C��(�7r��@�@�e�h������G�/�ă	����S�Zk��w�y���uݳ6�M%��LW�d����l��5�����9���*n��Bm�]O����)�ɶ��z������e������W���P�U�e3�iArS���kݭ���b��1��G^i�_;a�M������*5 xM� O ں!Z��~�
C}�du������y�ʳ��I����R��ld�)P���1e�Q��l2�n��p��\S*�g�l���N��*P��,���x2(�c���دd�k�idN�OO�^^�ԃy��g��7�"�`UrTw����	p<./�jV)���ʢ���&���\0���&VExW�����.���>,�����M��������⧭:�1��_����K��8��9��� Dk̽��x�f��E@���w�o�?�q�0 �������J3�]�v���~
M� l6R�P@��{������3��IK@�*����/B����#�����mS�B b�[L���xε�Ơ0���
���$�@lc��V�Ʊ{���	+�:��W�T����~�pr����� �?E�.h�-�ɪ�����(כ�h��(^���pt�Y�YPQ�i�Y���tZ8����~>M��������4�8����B`���*@ӆg!ǅ�w �kz�E3����b�����m�'����
d���Lb<%�؝I.�
�%౮����|��)-d�:.���Ϋ��4�X��L���?
H�|2P<E�BԠd�o�y%LK�� ����HI��M+ݢ�A5OZ��C&�H�D$���:��{O��qh�W��'����������l��e�'�j��L|8]q����m\]�%�nB������2�܃^��6J���Sy�S����F�69.�%D���,@��{8pP��Gc�A��up���1x�n�����m.�[��+�ݎ�7��K\}�$C���<�K=?w��D�=�Û%�w�xGI�[���]^�O9�U�#鞮��
����f��$/�����O���w^c�=��x�� �����'׍�i���QZ�2^f������pJ�3`�����X��G��y���0�Z��7FAA��V�0b�M�12�؉=�ѸʝQ��A�v�p���.��a{K��B�:�S��$�%9���n�� ����t�؅>�F!G���Ǐ��L�j��~�֣L�%b(5�9��{�={=��Z��y��-�;��t�lD�>}1�m�s�g]�K:.�6��' ���qo�|�0� ���]�;����\Z����f���}�BZ��#ܭ��]�#���=�?���!�\��½ʬy��ܘ���?���Pd��`��V�����/u�J�wiZD�'��nh]������b��*lN��F$@Z�n֢��t �X]R���]� �`#�Vkd\���>�I� �C����(f��D� 1A�6.��c���\"Cn	�|f�N����Y��J��K�4|�\�"*Ս�h��`�A����Y�J::���b�1����:�?�nWܯ�����R�ɗj�##2������DpѤD��V ȮE�C�-"�w�����O���'.�}g�D��~� %�O8l課:Tl/��{X�lF�ڡ9��%�[�Y�6���8Yĺ�4���.�(ԈH��5!�۫!�h���_������Cs^m�ذ'@�f�I�#�u�>Iw��H�'�]T �I��ÐCחx�gY����=�����?���u��%nh�6��q��2b��{����%/8����3�ߊ���Zuc�2W�
���yr7S �ѻ���޶E�����Y���<TցM ͈G����v]<�R�N�34���Fw*����	v
*&W��q2���b��l�s����c�_j�!�!�Zv�	��ZM�C�f�R &	�p�ڬU\�m����Wb!�l�Q�h|O8"����K	}���'06�#��5%0�%һ��hZ{�"2��&�3�H#�OX�tܼic�1řoH��qQ���u�-̣��a\@�Ъ�`��%v����*����A|���-[tiW�!C�﹕��v�Vu�I}M[���	�| ����x#덲)��( �1*�%�[�^��W�2�݊n���a���X��fA�a�F�~x�fЭEƇ�Nn+��kΘic8W��������)WSNlP�{��1L���4kٲt�\Z����A��T'P�H�J��V�.��Jw��C��7%Z�G#j9�����*Y`a�I26��G�k�����c>9�0\���g�c\���|�D�&��sGS�����{8��~��"S���W�z�v�B�_L�m'��
%]Ma�U �'u\�h3$)���kJ|�ءk�V"�B�E���>��5ub}8�XWU;����e�0iALIM�.��	e%��
��G[Tg�������Y	�1��B��&��PrF��}1����TJC=�C��	&�Hԏin�X%�j�[^/��߻�@81Y_׿.Dߧ'��/�����N��]k���?���T��ݶp�5�d��Ϧ�4���u�<]�G���ğ�n����{QHG�-Ø{����&�D�«	�MC�w��p	��8pF�ɝ��q%r�H�mY85�T��z<]D�"=	-�)�����".K�~ɰsJ-'@�kBe\J�"���#�x9�)�~-y�B��A�S����V�4�K���.��.�m�]s�4����L�J�rQ�DP�dHP���K}�*�M��HĖ���T ��>pB�uUI�Wr���J	���_�@�r�)u(٪��h;]O��+_��Vw,^9'�V����xG�5��NI[.��)�^��������	H-�1��ox�\|�����\��8�������T���"M�p�E��CJ(]a��4Y2�3�<�^(��Y�v�L���˹�n��z�?�?ːp�(�13���%�ʥ�if���*���{V���(۱���N���������;$����\�?��.�����Sh�/���(����P(ߣ�0*r�|e#�;�aĹ��ˠ�}���Z$̳ݟ��
M�V���L�_���6ҽU��W���SF�E�<���caƼy�����J�"a�?�H	* a:�!�	�}�ğ�/CD�ߣ�y=�t��A�%���{z�w©Db�ͭ��U!�*JNլ٣Ӧ�v���ܝ.(�n��\s�h[��֜�R�q{�]*��v�l�[��W����Z &b�N�83�w�5�`��e�m(^��Bt���0ؓ���Edت�`�3W�k7��now��, ��|_����"ҍ�a�ճ�\���Xw���Fa�XH��C�[9���'����s�1N*��2z���y��	͡�����bs�N층rh ��r8����ᕁFV�Z��Y84���ϕJ�����Ax���U�cp]�(Os�L˞k�;h�r�&���X�J_��_��+��ʍ1.�鎓/���q�N'�!Sk��9z��;���ò���,*W+-bn�H�7|^R�D��-��ټqW�ǳ�Yvi��� ���g���e�jv���2r�[O����<wu�]�Є��?�D�
������_�ݏ2��e�6t���Z��ʌw9W��X���xrJ�< �6�-q!ۈwlG�'�g*�^�I��|�t���-a1�sk�5���ֽ[��?9��ߠ���-:1�P��ϊ���y��A�����O9�$ܝw�א
��{��>W���5��y8.�}X�,��M����@*�?��dj�/=.』@�Y�,��h�j����TQ�1H�&,������������%v�".u�����5�8�L�����<a���
�k+O��a���8�٪$��Jd�Q*���lo_@3�de�u.M܇�k�Bt@�t���ꊸE��'��p��O\�l%���X^�4M�Xr��!�^R"����,h���Cȹ�aȮ��	�#����L��V�M=���Bz�����S����u@/"�׊���@�hg �4'����oH����%oi4����R0�+	&��j>j�.ʳ�Hp���������\M��z<֯";}ܶm���<O	��m�������;oezXbE��&�<.��.�Il�$D-��Ĳ0^e��d�)D2ʦ�>�r����j1��2��/�}v}둦eK�e�Ac�I�_�V�ӂ1>i�A,�84��Lt1ˡֱ-D�܀��M�M3����e���H���'�Cw'��^D|S��,LxM�F0�|_�4)���P����dABq2ݕ��$�1o��BIg���XW����A9s���έp��)lz��8Lˠ�� �ÌN\����s�߷�d�t�)cs�~�$���I�ϒ��Z;H�&��4ܬ��o<E=��� )�����c���*(/"8h������"
$�pK���ɪ��R����-��"�ϸ����SSi��V��4<_��,��P��`i�
gH�_� 1��"�(C�gb�(�IA�}椝��c8���[>O�n�x%`��v�u�c u�{����M),�[#M��e���� �քe�%�GI�m���v�;F ȫ2^��t=PL�\.Hy�Ýe���Q��i_縲^��X���(נ�r5$��GFL� ^��-��Ů-�1������	����I���T���E+j1�L-t�����9�� ����!�|�M��o~��$�QQ&fqEaJ��K=��q�G869�\��"Z���'�=Њ�q��i�1+b�̌�:�=��"\{��=ğ�fX"c>�� ;ڴ�c꾗be��\J�.t����H<���F3�����u��U�k��5�}��t���U��=�����j�XS����f�L��g��N�ϟy����I[�@T�4-Bot�3c������@�r�"����K~m�iQ�#��E���8寂�d�jA@öӥ�s��Y-j�b���;����������߿�=����Q'�q��,�6*���p�dx�=ە�
��wߕN��~��I���8�5��)%�F!�z��{)`Z�y"8������;>���/��]��N'q���h.�r]{Kq��E�L8v/��;u�r�^ �|�	����G�-���D�E=�2^,4<����<��7Zy��L(���5�8�B��ŀp�gF*�'�|-�����D.�&������}��,�>�^�`�UY�aI���4�"3¨=�\Ȓ��la�o(�M.0fn�Y[aRCB�h����:���*�9�¹����xEb6f|T h�v��ذw��MyI�$��
LK)���v���ܚ�E^(%�V�ΆQ�m�!��*�Q}�H�D'6�����>�p�Q�Q飣c?���B(�H��E��?�8�����]���oZ���Fo`���&.]K��K]T�b���p�Uz+�´���ƙ�z|㇯����Y偙�_s�21H�H�|��qW��J��&Ч�{E�*j�E63cQ� wJܴ ʩ�)�E:��V�ݚ�'Z�?)�{�1�j�U\ g�B��Eg~� �N[�&��jsV�&���