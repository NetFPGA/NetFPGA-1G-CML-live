XlxV64EB    7c4a    16f0�~���)�k�<���D!({�Bq��4��
K��;k1%=��W�-��ff���Ơ����Q�$��Hz�r=��'�r��/��}�G��E��D���->�-�~�~�M���us���03�^he2D���Ǽn�K�r������I.�5x�)S�
�ם:y�)�ޚ{R�ߺ�M�HB���ś���~�Gf�`"�g����M7:�����7�Q�팎y�x�sL�gц�5%��A��6^1��r�)i�ە3f�WL�1)��5��J+'0�����j����w��J�z�CFV7D�o� ��wӹ��?�=��.�L���,Hۨ4�����y�zh<rk@��O�#@H"�UW����~v[�>|����L~~��y%'5��K�bY��8�f�&?��8��[<k9��� ΍:�;w���-7��	4��^O�0�	�(��������R���{�Zx>�p.c����_��������>�tI	k%��v��k�o8e_vCs"a�I���.���Y�tko��ˍPp�0�4�TX�7H�@�nD�w��x{��j�_gQ�W�>�1#��[����wO#V��"��	D������k���ʱ�����\�&\��M�~��[�E���8:Ya,��܀�m3�[���eY:��T�®�<0�*k�c��֧�ﰾ�N����j�v��g�&nQ?���km���૵Y�|l`�)"�)�J�zXb£9?n�b� ����o��T���(v���wd�!;���N����rhW^�n߆�kY��jH�3�	��2����亯2(��6�#*H���Y� ����eJ"�­DmX�$t�zH!G���{�U�d�2�G;�=��h�������>��:�:�1)�<4b�+���B�ߙ���>� �E��8G��ϒ{���\y��%F��<^X����?�_\�_E��"ό�k�n���j��\Aɽ�e� �GŞ�a���u,"���0Ep�|FLj��Ne�]�B���&@�ܡJ�֬ӟ�w�c���0�9������1� k���j�j��d
�z,����d��;�v�B�����Ċ�^��qr��X�tF)hwF���rӶ����xik���,@Yj�ʍ�T��=��Z��	�2,�{��l�.9]�Q��� ^]_�l��"�EBp�W��;�����8)8&+>5���}k��R��$����"D֖���?" ��d�`�`�'p�!"�E����TB ��?��36ǹm?�"������9�_�)�3�#�>��g`��l=��ȵ˻����p!��mnXx�Á"�L�2��%!,^HYy��T��5Y*��@���)��<)�I�O|k;��]�p�v
y���b(�L�v.94��nUo)�1
K�JRf<PI���A�Mu�|�ym7P.ḛN���X�����	s۪�d�G���e?6�m�E/���-`�����P�S�x�_���4g�(/8�J����(Z]�5��j� �n��A�&��9+�b0�1~:G\ꑈ��Z��Ҋ>���nt�4�\�z��]�g��Z[Vg��[*�s�w9(�MF\V�Z�ԡ&㭔�Z�K�eg����;�/;2�O|��Ym�0B�"ޢ$;N��N�wZ�3���S"Ṓ�i#X�,��͓Z��Is�����%�"i~��������#0!��G �u�W�ē��e	�y�B�]��q�O�N8��2�ʿ.Q�#��%>ǩpf�8��:g���IP@�"yI�y-D	؛�|��su����ƈGy�Cy��A4�
�oZl�4K� uCo��xČ���ٖU��]�ǣ͑,�	���P������G�h���}uh_�*3N�Ku�|W���;�K�����~*�=!To� ����uh�dR���;4�K>A�b/���S*VM�"�������3KEKY��v8q�U�s���yƑ�aE ?���ЌЕ�2⌋��E͒�ߥ��Wdq2X��h&���T������l�Eސ\��i�Lf�&�M={\��Ѝ�_��zB䴆�\U)M�A��	D�ՙ���:��HH�,�tr�P�A�x�h�6���}W3@��7�аƘ��g]b�j�k�tE��>���l��wp�y�;�E��'	�	U90�4^&˳Sa��sѓ�ܣ�6Xi�^a>esk�f|��)5�X[��;Ǣ��)�~s�	m-�Fp�x`x�x&�.=� [�&�F�o��RI��}����x86��P��}��H�����#&�T��ֈ�*/H0�e��i�;9Vc����Q^�Yx�B���'f��4F���y��7R>ʎ�\Pf��%�Y�L���*{B�t�E�ڠ슊W	�"8h�����B���S���O���y2�ؖ�AM�S9�O�G��
�?�LK��S���~z&��_x�`�<��~�|6dʬǈ�K_*O�ձ�ʓ���Ӥ�Hȳ�04[�5��WE��P��5h��<����9�G7�c��L��9f��Zt���s?.+x�P�g��(�ɍ}�,X
���@55{��`����K��L�8{4Ew�4�T"� ,Xz̓�	Ό]�[�� �^�l���0��ToRegftQ�� 0�"�vC��&�kb*>i�^t�9f|
O��BEr�d�����A�/���ee��#��K3�]V��H�t�I{��2�}"}u}�k:��P�Q2��Qv���><�.��#�����R��F���O���Pw�R�"�O�9i�(zx�j�} �E� ������+�i[�۞�<����	�C0�pv�S��^�cO��Ї�!�TX��vl��l��۫kCt��z��1�*0���v�,����-J�hԈfϻ�A�I�F����¡��!�
�:%�ku�l J�Nik��v5ȅ�����VM#�n��}�� =]�M|%R�Q��w�3�5�B���>?%f�C^L�.��8f��<;�$Wcd��n�KW�A�P��*�����v*�`8��m�~��k�����u��|J5_�߈8|Nt͞R��㧨��,�}��k�:y�-� 	Lv.e}^m�t5�lF��3��J���v�����%�Uⴐ����������(R�VV���%(�*���w���'ʹ�����"�i��&�yт���)�>�6y"\�X�>AYam��ѬLa�%P��gӻ���BT�z�!��%��Nt�mJ� N�DB{c*�sPqKt{4���ǎ�|��]hCQG�z,�C�fZ7N��ezmR�~c�^������_!�q�.e+���"����;h� ]Y���w+���T�#hn*Yq� �8���� ǜ*���2C��'z�=f��c��j�P�_��L�l ���xt`�4)�����_�V�x��K+�??u}�����a
��i:��YE�,7��s��3=z��'7��3i���=��iii8���̽�Y&����P[/v��>�Z������b]f���h0��x�V�ؒ@%�ƻ�7�����'|䵶�}!?�m�fT
9���ґ$6I�U�f��Гˢw&�}�Z�^k��o}ç]���`�]@hbA�\n�R�f<��.��)���v� ���z�/R��fJL�h���u5ŉ3檮C��+��,�=#����˶���t�e�YN>ݿM��!�j-�)�T��&RdDvҏ#z�n�J�r@�Z���P�c��M�,�4�8��G�
�
��cA��C]���ӝ�(!�5,V7 \8%/���=��r�p�
z��C�LB(݋O0"n�g)���U���?�i%J2we,z���F%��DBq�r����L�<�<;'�U_�I
�P��Y}2��MD�ݼi0�E�ݰ�Qf?p�o��>	9C�_8ڼ�$+�U�8.sLuØE�ϓ�z�6�����Nh��K��Yq��e!>Nr����F9]�D��[�������S�N�m��|/E'	��)���f�kp̀�s�X5�g��7;�~H���?�̦!o�D^Q|�_��������|�������˶K?��VDg�v�*Vw-���D?ZlEU��0������H���hȸ����MT	/��>��-�����`�C2�!��nnW�}�{-��{�ª'&�hw�RѠm#@CK"dF�!V�Y͗�;�f~a�|�߱C��})d`ә5��<�W�h�����&
/����x�H/�a���@�x�E"�5�]��!���Hx "��*�Q�j�*�=��F�?��D� �Z��7��C�#�.B������\L����R���&= �vj�l��ť��B,<_�M�S"�3B��%k�-�-�K�k�5���w��v�PPv���m_���T��RF|Bo��z� ځq��^�&���l�1����k��!��F��=��snKU1�J�{�̢��~��K��1S��P�ͻ�B��L�6|}�Hq_׺�tޚ纾
 �4z5u� ��~��C�s�� �@8˾�����紓G8�C���
�;�N��؄+>�+kn��Mk��S���cSwmΜ��b����-x��Q�B`�|aoc�
D�Ei=���%��&�M`l�ԬVw��ޔ�f���Skg�d5�=����!,�԰4�:�X�	�*j2`��E��8܁� �����w��_b�ӱ�LA�ߎoPõ�̲KA�wq]�j�g@���̲̹�X-3:y�*�t�%>��B[|�j�lI�"J;�z��|��i�o��8<��d���Ag�:�k����Zs]=N�iTl��=m�n��D�9�q�j�bjh�v���M����Cn ��������6�6���A��P���]�/ʀ1�g��<dޙKp6w�����$�����ąf�%t�:e����Q/y��Z��u��~���lr!��d���|�;�_�!>��n:�F/��c�&d��t� h��T���dq��)��E���xI�7 �zC�O�6�xO�9�D�0���������;����cB�N�X��N�.���1W�h ���|S���<��˖r�M���G��Xc �7��P��(;r�Pj�&�:��Tu��Zh�/��6��]��~2�s��#��q��v)Ȩ��(ѵ�1{v���(&"�͠z�#��ޝ�U]?���@�ťO�_�0�z7:����veru#��bm�OC�$a��s�+�m�������)����cO�;Bg����I�JKfE���ƕ�����۹4�mL(X@�W��C��!s/r�Gl��8˨k*7����K�N��ƚa<�1�86k���v"����5F�g0�
���;m��wJ���?�hR��*n��㡀��n�:�k��]�L: 5�"q�����������Û���ZkM��m� J���\C�hɐ]Ù.��@�؁%CZK���p��y��$���/q�d�}ҀJ���D��<��ьR�5������ؙ5�Bh�lۢ�dR����,�oc�9Nw�G�p@cuּ�D��`œ���ow�"�S7���E�#2
%c3�z���HC<m/㕌܃��U4�Yf�&�KN�<�V�a��{��o�o<>7���.U^M�i{Ϸ5�p��[�hU~��w�07��ݜe��q2:�z�g�k3��c�~@����E"�k�;����#~�Sˊ�����E��9�	�"��2�3Y�Z'{�!z��Md��$�~k��5^�!p�$�~��������"��v�1�F��;ϣR�l�qsR�OXO׸��3�a)�BO�z,Bm\�O�O�VH��rEx�O�0�}�`��$W��N n=\��1W�Mn�`