XlxV64EB    c9d8    1a502���:�*�\�W	�p������1�����U$���������S�E]yKji�A�\7fu|[�g1�u��ji�\��0�2�߄���T"ʙ���p��K�N��	h��]�w.2��@+ο�U�L;��ʲu���5P�*��N76��y ��I�o�t���0�T�c�K�6u8�����s��3辣x2߃�CV����zr��I`���԰�G.c? ���c�`�>�.nm��<�h�tB���+wB/)cI_`�����}'�o{(�W�@<�D��U_nw�Lq�� h|}����,��˂Рm�bG�U�y|�!�N��Pךt9�{+����3��P/�1=uPHq�� 2Ԝ?�$��Ej{��uR���@��(�Xh������d�����qj�I�<ӌ��T&g
2� ��J���>�$zl���!��� Z�0�ة:L[)O@����=q;Hf@16%:���o��Qu=$���.����0&]��A��s�W���bu�
� �����/5��f�x������ŢlkU	��>�IV�31�|�)Ru��ǁf�S��*1[���:0�~���D�i`ݎ��

��r��eO�g�y����)"�m:��E	�&ʔ�=};M�U�<m��2�l/q��c�֍jZ�.�Dٵ}݉�LJ������̥mݝ����zEH��] A.�w���� &4nI��׈�'(���A^��c�b���zһ��<C@]��&��1ӪO�S��F���~-�6y0�jw��I�^
d������B��8�)]��(gL	�i�&L�LI��q��Z璕�\�)���b��*���5E%��$���gi
�B���c#$��ե|��f�[U�q��7�Y���s5���)�QG�1Z'{_c4�ۋOo�-y�L�����=I[�#ʆ}��p�s�A�E�M�5/�u����a��+c�X�@L��:ZC{�_���F��5�Ra�i���V
�f�Eߝ�-98`H*jN�B���	������_�2� S8Kk�A]Ȼ�y��]��?�N�h[6�>���ݱ�%�Tge7\�HE/Bp�sz�:��CL4����䏽-�s����4,w8�l�]�M��2G	�k/��b��sߚ�S8�	�/��W�sn[Ū�9��Pt�yP���K�V�_�6k��Cba-��A�s�
�m ��&����7H:1���lsA�Rt���ϮPp|a���Yf;����N�)�Ȩì�b�Iu�R���6)�"�u����S\jT�[�n��������ʋ���D����G�>w����fpȃ^vT�+FျO�E�PC�/�\^�g��su?�P�x(y���� �������/�'��z��)�oY��|�O�/X�W#Yì���cZ{!�$��b8��~�j�N�܂؄�ƫ�JRrPC�m���C�`�b1�N�>j�̒C���>
N($�i�\��L�t(��n�+r�]uN�d�ug^�5��S�*����݉i�Zl�������S��ޢ{Y�uT�]��t.p7�� ��?5�<-��GXZ
(�(\�/�� ]I�6�|u��M�uj�#a~��<��qn�~Q ��}^���z%����i����%J�4��췃ޜ����\DGpaFǀ����M2����aϻX�h^x�h?xȗ�����V�Qg��H:{FW��"�Sk�Lz7D>1J�[1�.Y�`�ۅ�C;�蹧K��TǶ����8{xI� ·R��D���nЧh��E�RU�ۍ��k��gEX��L����$�{������u~�Z��n묍x���V/��
����</�:�R��B�N��~,΀�!� �)������`h���K�4�*���<N�1�CwV�v��Od���Q���=����ٟKw�u���9�h-#�ɷ��`(�W��"^La�I���7�1x5Z��ك��l�O�L=6b�I���<���U6뀊?k+�M��e��:�"0c� �ιc�/S4l�R��Tyrm�Z��R
63X���L4�~�?u�o��Eo{�����fO��6�֝��w]�g�x��p��΄�fν'�e�jНúz��f���G{l�Dcj��R>������3�=f|��9�,a�����'Y r�7����_�%r��o��Dr8ׇ%�@H3X�0�?8(�/�/����$M�n���{�{C� b��a�Gܪ�2�-���<��z��"7�ø#~	Hyn�x>J`D.�$���G�����/��0P|�o��_�/kc!�q>@�����L������$�w��f0��ݽ.X.�xț�{R��_����x&7F�$��i�&��Ӝ�� f��Pp�C���[s����F#Y�R���ȿ2��h��[��.��z����<x:|�`���t/�	�0�@%��E�R�R�W^i�N��R|���
Ղ+�<���AK#����i(*�?�ğ@�E!{�^ ;i8A��a����d��<��N0���'pg,���1P�q���Ab���N��d<kL��p#�3���ۋ��\��P��f����t����x1���GIŲ/@,���Nqbqë�W�� Y�}&+���>�,Y���*@�im�,V5@��rr`��u�x]�؇Cǎ�\�����[�`��MէQr9��׳l�ך�G</��SQk�^|V޵{}	��@���� .��$��O������j��7}�����h�� ��>���4�T��%{�9[ �"��}��w��ڧ0�S+:�4&��(&�Y���0&�h�u�@DS�6N�Rڸ�t(_<��ס��V�*�y7>�:��� }�f�.Մ_��uc����5C2�Y�s pӾՇD�����\�쎡�En���A&�Xip.d�ޮpk����{��ox���q{��O��۰<(:��o��"���V%	�����Fz��`�x�fd)�AQѭ��h��y&MlFh������|$��s*"�+�aE��밮�ô�Z��	�Ԥ_��M��i�6��H��'̽$+"�"='��,��*_��K�[G�~u{ɞO=RVKH5�s���5ǋKJQ�@5i�.�V����|��c��'���<X1�d��a_���Kۮ��MI��Y���,��p6�u;lJ���ĸ<$�^�j��8��0�TE�Y�i��l����$T&�~�xL��E66��*M_ ��J$�hp�R��=���{�]#�km��c9)v��4�؉K�,ۛ���%<���4$��?`NB�]�A93����ܐ;��q�S��q�J�U`��8�ݷgޔ�D���V�k�+bW��v=ו�x��Ng�	�%P�9���٬e�p-F�i�V�@�}O�x��k�b�ɬ�)�pȞ�E16K��Rڮi�R~0u�Ӏ9*I失���j����S����8LO�X^�3)���y��������p�^+_EZ9���s��}3����݂��{��ۿWd��Z`F�*���h��+�qY�I*�$ۊ�r U�?4�M����ܨy��n�Gs_.S�%V���d*�;爧���:��*F-�~����%$l+�p��i-���`<��Ƿn���� ʮŪ��'�KP�z�R}Q����bp8R������0�e�k����iWQ$M�]�iC��2�R��	��'�·�����siۇ��	�E�a=s��n��� X��A���ޞ��4@��u���:
\#z8z� Fr�?��h{ȑ"j0Z#�ą����1�ǐjo*&F��YFaXx��}�*�s�}�Z�	��0�{Em���������81���lr���$�ǵ^N���e���`'<s�ZPZſt��s�/�Ts���E�g�1xفcO��)Ǭe Y�6{��WX㱊�#<�&���S�:�oKd��������W_���,����E��^�%�y�y�����+�®�w��f��XXI��S�fj��Jt�Ts$�o�5����\�C��@����ؗ+n��|�jg�o�x�R7�7�Ș��#�ߪ/kcW7�6�E �#D�g�eB*��g��>!$
~�@�<B�/�@/ɱ����x*B't��eb�&��x���}?�N9X� �Qwӈ��3HQ�+��bQ�2��U����a<�" �\� ڽ�^���j��~�rD��-��@$r��n!��;!���Yp>�H<��2Ⴞ����zF�������������5���RmNJ�d{��x	ʇz��hK �sFu
�y�TF��˪`��}�G�&[�%�ң9�S
�]�Ux�i�0{�A�7Mc�G���h<�>���f';	�{i��<S_����F�@HQ���<|p� [��T �<����z����&����$jߥ��R"��Q5]CXD6�O���ө4W��9��ўPiD�w�0�c�Z����5�^���Vu���0ş�=ٗ,\�"&"����L�|<������eY�?��ш�ɓ��>է?q�$��O��Rv� ��➕A降�O��J*�򁵲��<
{	x�N�xX -��0�nu�9=	�Be��=�l�D1�-����v�ϯ��i��ְݡ��c2�9S>��`K�'��'��s���ʿg������Q�Zh��nn�}�����K�݉>R�'R�*��i:�BB"Y�N�S��U�eACXz5n�xQo��y��7S.�Z_�9����� �u],���M �'�Z��(%�>k��p�9�?���܆
E�r����͠�U|�a�=�M��r:���f�(�Qg����}��!�U?���P9�4k���J\�	T�ap�$Oo5!��8���~ho��~]Uue�SN��^��JU4ճ�W�T�u��G�1���Ń���(�Q��V !<����x8�Jj��X���-�g��T������VNo0��Ss��F�5�}�@Z!���4�dJ�0�RAȲ3�\MXU�ٸN�ayz_`S��;<v�Ve��	������T.�e� ����b`&-m[���Y�賖DetWM���TR�O�Ee �<hP��~R�f2ɚ���=�Eb6�l��$����ZM�iN��i��r��u�Ex��(3�gkU��"4u0�w��`�m_�$���hŐtT,�����`S������&va�S�M��h|��L��
�W��ę2/��
l)��{�|�Lإp��m�,"��tI�\�\�O��[��n��#�xI��?\������[�Z��$C{C��C�3�@\�+��~c�*����� ���L�U�Y*2n,���ny���}��@ �M[�rXݏ�迣ֳ:�!ӣ`E�!i��]yMXo��)I+���D���$V��|G��1v��ʢ_i�U�GA��p�Q����(�`�J��� �e;���2���ۯ�0�$FЗX�)U�a��,V 	1���7XE2v�\ *�K�?����O�1�
X��8"�p�G�v���erQ���d�ZF
?+�[�������u�jn��W6����]��&g}^����
�s��sC���.v�(6�����`ɺ~����5D�[�x����9�)�Ɍ`FD#��n|�G*���C)�!0�з����
�=��S��N����8��
��q��j�BB�l���-�pzu<�AOZGQ�H9��/��!k�E-_�ں�� ����K:=�"2����$�x�r�ܮ�6]O���k6�/H33P������eF�`.���X�JS�Wy�C>���3������s�Q��c��w�5G�y	K��=�X����ξ��=�E��Z�<���h�P�J>��i `F|�a�*�� ��ݽI^7`.��wٟ
��^)�T��̘kj��M��G<&AW�S0!0���+.�s1HfkKZ��3�X�؏P���EK��0�L�D��"\��.)��x&����u�L�ԥ��MNA�:$�AJ����,��
�!l�5�����#�3��[�$���_t�i�aR�|��ڴ/b�9�(ގ�nk��3��P�2#j���vު�~;�Q&��q�I�&�2�W�Y��2��[��M��F�O$�<̧?�+�[*ʚ����fRJ3��' ���&BQs�x��i7p_�c�몏��W�Ν����z�7�����|٦o�
r�S�X��u�-��ƣ������&��M	��n��u���{��#Qx����N�#A܍,�A��CpE}�s�Z���i��z��F��e���$�J�Oj����|~&�~1�b�[�~��y}5�]!�F�:��hV|���h��l|����B�Qv��GU��a��o2Z�����;��f�;Ȕ�=����I�J��I2J��q�?���ӹ�O�@��,�$���%�f�����ƄN�@�D��[�R��C��Ҧ{�0�� ;�jT�	�.u� I����䅄�U�d�c��)eI��AR��䤢�&o9�f��Z����+����XE���Cg
*k����d��6s�����%��5��tt��r�c-_w���A��F嫟��o(٣|�x:��78��a_K�LC<�[N`���ǜVS�!WC�Ÿ��	��