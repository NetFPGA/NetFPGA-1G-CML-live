XlxV64EB    fa00    2ef0[w��[��rr,���;�zˈevd��`���O(���4-9a��M����E�t�M��]�&���wب'Mtnk�9�	���!�;�Y���p�I��R�O���W;��0="�9!�I�G>i?w���	��9��wx1�G���L�N�zE�,7w^���R^��}O �~}u���0�Ó�*S��p.[L�ߧ5`�n��5����`�nyE��� ����[�9��q׺��R�@�7f��e���A�O:�2&Bt�$8 _CW(�E6��̢=���_�>�P�9�c���r
��Q���#-&CM�W9o�p�nv:�C�J��P�X'6D#�C+������$�l����v��$#~�f���0����vP�!��M����@��f@����<���A�l��rM,i�`S���5{��ԵO#q.n�[�V�T��4gB�����|��ʝ
�[�:�
zw#ri��d�z��mI���<�����]#Q�o2N�$>�o6��$�N�j���A��R�[����S/�_ NI�D����8��A�p;&����KE��^������
 JQ���� O�4�~f��hT��_�_�zav ���[՝�(�� s��e��S6*�X�*���fF�bX{2��
T��	>`��ȁK��'�_n����B.o���L���	�aÄ��{q��nO|��؂��ٜ�G᪏�:��
��3W�Ie_����T�_c���#�B�b���R:�&yF�°�N*Z���'�� �$jο��ר����o��a�����`�!�d����L�A���;7`�?{f�hsq�,�0�0��&&;Q(ڡ��j:zڛ����f�,�*d�u�o�1�.d���\�̕��u4UH��V�	��oĲN ����o +x�/���Y.`_��d�!^�T���gpm��\�� ��FqQ��d ̅��*��{9貊��^O*so����@�>!nUg���5f�E���P�I��c3��Gt���֚Q��hS�+�����i>:͹\GrxWb�n=7��g�f'h<Z�)����S�*�YX�YP�����a���2[��-�H�g
�Ĝ��a�9[�!Ԋ�0�.좶3M�,X&��i]q!�_1�6�x$l2@���c�I�b����<��*�ڂ�u(L�'���`LU�0�?��š�?�Izg��D�G��ݴ@$΄z�#Yw�o�ե N�s��m�������R�!0�����ӫ;����w��r�p���
 P∷�]`��Ez_�Iо%�� ���.HXv�����Og;x� ⺖X�
���3h�O2vh�\�mC%�������0������%V�k��@��ԳŔ�ƻ*�:d�`l�V:�����"[Ű^���[�e|��r����ya���G�C�w�}���1&�'>!;�SRf��F���� �L;�`%�xI"0��K�cPN��~�&c冒�29{���g�0B�;Ua���bbi�B����ꉷ��L ���v]ںTR���-�y����ԓo��8�t�yJ�pܪ��3��>����$=Z��c������[n�B�^���U��<U~�ڣ�Hz�a���o ���s4j��h���!�O�yQ8Ϯ�^�o�f�;��I�Z�ź��gF�в9C���K`�rKW5-��|N�n�Q�����,�dL�!��ޖY.J+l�8�XK�����:�5����Ǻ#"��J�O��2��^WE�ǉJ�ސ]/���UV��EO����)P��͍,��O�g������d@��y�󬷵�ʽ���EU]����\D������S�+C2����GC:���&�!s��<�T�/[{d������ʚ5R��r�rІ����Ut�&�
l	V�5�$��y�5�^$��GN�r�� �Pk�ל���X%�ŕ9��C��ꧽ�U�r7D�F�[Y�7��}�5k��Aژ�<��y�6d�Wb��K�<�(nc��:yb5�RTM/�G>�>���a�^%P�BBpS��l'-	��� b�X�$�����ݘh�D��KE�fR�|���>�A�^�B�Z"||��pM��O�X�ɠY�uADAH~�.^J�??Mq��i���K�nB�NvH'����r�T7c,q?����r2t�)�H��L%U�4p�R� ���D�v�����}љ��i�МW�����L�츹�].��6��A��KDfQi�[,MɃ���$��'��¢Y�@+Hg)n�?T[�M��F.mv6K��:��p ue���=��w[�����p=���x�q{S�Q��Pb���f��7���a�?`�|�|��M� �.�֕��UG�/�c�]�t��v�9zk���Z�{ϒ�sF�ߔ�����ã<�9���\ϧ7U� 0[��VǛ8�[��|E��h��������.�_�5��
[~�c�wS��m!Xo���n����r��,�$�@u�b�Ѷ��xG���U�҇��)�oi%�1S�	���"F���~�%G;��`��5�&��z�U���S����A7�V�|�y��tK�wb ��u�k�M�� [Zy�IWG!�D�5�=�d���r�[����z{�+"y��V�d�_I�$I`�� �I  r$G�g��kڛj��+��F�lG�ʉI���;\֗�J�H /G��#V��$�M��\�['K�����u�@�4;���e,f2(���&��u�m�i-���E
f�SȎ����9$����������q�T{]X]����d��JNf�[T�x���|�v�$�x�_'��#DXf@�m~�t�f�|�>H��6���j��R�t�I'xLp���~�n�Dm�H���.�bƍ�����ǮqG��f3��wx�'�7�	�0L����x;�{���',��r�� H�"��Q���ؐ�������4�s��M_���s�{O�XߒT��d8�̸��K���5v� 3��Q!F2A�̊5��T�%qU$�b�A�a�b��<t�DcM���܍x�6��FQ�mB+���0�a~+vj����uX佌�/E�i:��N<q뾹���X��c�ߥZ�B��|?�	�Od���Mަk�@z'�1�y�+u���%L�ʩ4�M�&����7 "�*�S����g<�x�����D�ys�FX2ӤG:Ӹ��db ���U����QO0i�Q�/<[�5����������[KǼ>�0�X
����~ͮNT�`���������~`]ɧ��weU�h ��[�2*R�?�����~-|��ts���D�\�KR��W�x�'�퇆��E���ck>f ���R}��E���h�S5}�s�Y)���-R�}.��֫���Ҿ�A(���Pe�;���Y�8�'�b7�q�9�=��Ai�F�;�gS|��Έ3)c�ߖe0�O��!!�7�p��D���� �[[��d,�;]�/�`?��0,�/8�Qd4q���J7J��u72I�;ڣ��z�w#l�W�x��"2-S�q�;b��#Rݲ�����:�W
��s0h�iD8�pD��:��	�3����LL��<�\�Z;�v�b�Po�2��f��Z_'�R���� ����M��N��·S�E)�T�Ĉ��H]��C�Q@y� "u�D|��^���CT��%��W�1���2d3��%�GÌw�G.����I�X��4����g�����ؚ�u�F]S�s�K\��7W��V�Z2��>�#v���y�4�W���m���o`�K�N���[s�F�M��!�j�	�O��fٱ���gP�����a�ޛ��i�����Y�O�+rŐKR?aHU��vo��ʼ����i�E���EPh��O=�8�n{ح�(F�3�o�8��V�p]:�X�S��k-p��	���⅕V:\��9�\��>:����7�3~vL��=�b!�c�gg�np �h��X7Z��h�H��`<����:������S?��
�Q�b��.#	�B]�i����2�t�?.	?�2���S���Z�:��>@�F%�Xd�;���d����o��vt��)�)�}z;��x�Y����t\��3���J��oԗF��{��j������ݒP�V�9�¥n��ɭ?78��F��o����@�:W����!U��ܗ��t��~�<���K�&���m'�>������/X�.
�	MU���T���[��� Lm�|�NWgۯɥ��3�O��h����K�0��;�rx�}��^�`0W��ī�ί_8 (���ࡣ�/q��� ���]&�N��e�q=���ðC��u�z�	���?��ő�k鏰�&�j����Q���QKG��eK����,�ϘBf����=���~M�f��ꧠhi�If)���K��s��?��B�i��>S��lc���氵�gx��N��!Y�
ö�N���m:�_:!p��C9�u�]�d����3T�a�14]�vWz+�o�٥+���� ~�$>��j�����������p�؄��9�3�w��\��u`K�c�yGD��P����k�����Ӧ�g*lTk�`�����#6m׿�>s�B�_:�{'�"f����� �K%����^�F�M��i�ﲨA��~��W�ɟ�Ѝ���Jh�1
����hZp�ڱIJ�,��)�G>���'Զ+��GΈ � ����5^�TP֏���	ɛ�N`|ث,�ȥ;��8*�x<���j^��]ü��v�E���W���X��g���VYqg�=�4d��̈́�B����H�Ό"�r I}���о6�x�3'ιpB2��$���"��u�`ݑ/N�)+�3���gj�{l�| ��H�7�N���7l	e�q�*��0��@���P�"��>���n��B�<�V�5�#?����GE[��ZyV���#ԚΏ���D��R�'V�$�}�b]|Ɏ�\QV�؏��w;~���!�G��/�h����Q�F�#F���F��V�Z�=��a�w* E���s�W	<�DiX��l�ۻ�Uuo����zmmn��X����=�9&�=_&�B��|�l�A�+f�Q�y�6cM�F�7���i1����FvG>;�մ=:,�([6��
����M}m���|�B����`-GŖ)�
��*�U�nBe0e5g'QK%(���]^�>M4Q�+�#3�;��١�/6���.b�C �}��p@����h�mz����~���Z��ծuanI�ٟ�.E8��׶��aR�|I<�{+KK�v}G�wX�_��sL�Oe�Gb�p�L��4�
_��J�$m��c0C�l@M��DP|$��^͒�=0xۿm[]Tx���w���B7S�3��Ϙ� ���1��H$H�$�qJm��+v/��k�!�!��Ὗ�Σ��Jx�R;�#�t��y�Y�=��CB���
��T��|�'�Is���_�3���HD���d�fⳕ�\C��������b\8�i�n'�?e�G������J���w2(dU9�����J�p��TK�w#��*�^y��@�H؛�=]i��	��{M��l>;E��>e�m[z�t��sM�TqFw��[��0b]�rx�C1�qv�Ru�*�b������J����f� ���]��J�Yfޕ���O|�	�7&$�,z�r^�R*�.�cQ�|����)�q�M�؞ir��F�_����#نB�^�:��*�ozS;�����n#���8�G���B2#Q~88d�>�;!�HS1@9��(��^C��+\m?�e&�!�M8sĦNK�g}�ͬ��o �j��Ҿ�E���Z�ş�ŏnP�C֟
�d�GS:����LH��͂�?���@�>
9��z=�{��}?6b��6���Ӽ�����|���v�0p8*X�o�&2Yk	�����0��w�~�QH1�_�B>�V����ɘJ[��H� �L�R�ƽ��ʸlї�wB
̋��V�� ���;�ʋ�XK���\��c�;�L�L�/P��"�Ub�?;"�V����z�Ħ�2˭��卓5\���u�(+�f�]yW)����f-s�Ep�-���=y�F$�NN�x�ZƯ���1<�� IB��㰅	L�sX$8��.T}CY�N/�����)�.��{Þ���NIJi<wK�,Q%���E�N�6��eH���C�3~�(*=sCz5�Wzm���p-b�W�8�B� e�%-
J�Y��F�u�s6Ts���@���+Dz
I�%�M��?�. �Ӎ� l1n��)�<�k��X��4�%��r�U]f��/^�'���Z� b}��)��]�ƜF���V�W`ɥi�z@2J!�SoS�֮cD��C

�+����`��?<��R�(��c����i'W���j��<9r%)�����.�W�������M���f���3���B�}ȄT0����0�����x�dU����؀��� p�Xǁ�ѧqv���Q���ݹZZ�$��Ҍ{=��d�B���P/�n)��e����:���u�ㅏ�E�[��WVض���ύ�_$�C���wM��9Q�����^A�M���OgY�MP��]��%�&tj<y�(6�a@,J�g��������J<�?\a<YD�����+��r�]5�( RG0U�����ė�~<�j6��v�F�Ȗ�z�ь�W�>b)�;�~��O�Zx�rJ����D�F���nQ�槀5϶��cFË�{ݤ���J_�;��=i���x�œq�v���	0i����r,�C"4�\��]�t�����ۆ���B�xZ�2^��lYϿs���iT������3_ߴ�TTf��2���a���kQͩa��&���Bwp�lY+�J�(!��;�^d��b��bJMB?`�	ӇF�r�	 �TE|������&��'6w�Ab���m�������+�o� 
�r�"


mD�����ޜN�ߏɅ�Ĳ�Ǆ�2;m��>PL��X�S����VN�f���e�5QKzGOe�f�$��79'��a��-(��,�*a3����k��^a�Z�Lv$���'T{u���F@mi�-J�u��#u��2�(����P;��0�`	^a�����댹lf[�K1�VPu��CiL�L� �u�����W&��B%a�!1J�q��|f"��!�-�#[��ZF{,?e�u��yr�Y.�%H�4>�J���)C�y�tظO����!$�HI�&��:Y�hw��hì�-ն>��u����jP�k-�E%e�����Wv�5�3���di#�bP�/��$;�E�z�Wq���g�hϚ�����;��QPe���rx3}�/��-�\��vԺ�e�A���3O��&>�`�`U���I�6�QU�:���=�;.�R G�d��\�r�k�Y�g�U��	������ޚ���}������x�2�'Xl8�+LôԔ�|�����FU&�����wB��`"��5�H��$�-p�9�9�wh�ީI�>����@���v2?��r��YdIX�(������u��#�&��˨�u���B��Y��傑G���C�����
�r_�N�p��r��SnJI�^51#��hú�<U:H�7?�߀*�'�v9���d��+�%!H�E:-�>1�U�\�\wB�юɔe� ��o/��7�	���]����\���	!{�G�8/_w��"gH� �X(�kP���%��Tq�٨|.�]��K�����
i�cp��<���n�V�P�,���բd̡i�!1t&�� �5 ��х��j�u��(뇾���r��O�V.+b�4�Y����nh�D���5�:l���H��#�K~������)��'��`<��"�q������I���|p��NW���2�#�z��2o��7mb�z���P�A*u�v��cz���A�Ev��Ea�f��N��܅�Xu�Ř���I���4dr���m�A=��W����x����IM�G�:Ԁ�<"��V���񝁙1�/�);
&����S�<Ib���6x�����-�v<�P�(��i61/mI�߹Tn,i&�08�W�>_�E܌�!�ɠɠ3;�vW�R�a�	��H4�R���a¬{�5�E�$����?�"���@�ĸ6m����,H� ���Zp�2! �iw��}�>w�G��/����[�b�8���ee�q�'�W�������8>M\@�v(���mM{o�ŋ��ڱ�<��C�WӉa �h�
n��Ӊ'*�jDo�Uv���������r���>��upN�C���~�ɱ�'*��_�-|-~���Ic�u����!�g�|"�7�1NS&�"l��V�Q��H~C�/;b��=r���������Y�(�X�dЩX�]����3���x='����k$sUu����ߗ��3�L�B^:&'/+�~C�S*N0�љmt�("�;�$�B���ה z��oԾ����r~����qZ�����������x������MB߳0��+�*#0t�N���#,�	HV/���6v[�x���l�%��'ʞ}��vi�@�f�#����|m�W�Т8ۢw��F;���As�!ʭ��Ba������6���c�t���)�m��x�-az�}��c�̅���|���B��Z���P���*Q ǂ���æ/*:���q��ib ��tm9h~����R� nbgM�N;�c��1!U�B38t:B���?����H��]�sd��z�){�P�x�ym��n	�s��ϟ\Ff��ZR|*�������g9�%�]�#���l�2Ե�字��M��;K4�
�6p��;	-ސIiP�˽\���W�sn�J@%C��M��r�Q���{�P1� ��wP|i��9ֱ��^��xҽ^\*,5�P�>�2���L���4�`9c���N��|)+����sU�c�!�_��%~��.�R���%���=U�P�+/��QB�_��-����r,�fu����0���_�,��ތ]����?�fu>J��� o �G��H��2��bӫ�����oص��$�-�I�Zw�b
����~��f~hq殣��]�t�!�gº��mG�ey�(���|��u��:�^����+�c�X�*����1~�o}9:}����Z�.=����g��\E����ޥk��-����wf��-'�T
���_�,��D��7P�RF)��6�$��ۚ��
b.�]��:w4����4�4\�`���r,� R�s�y���S���̀�ʘ?�� ��cQ$���^$ �˅}�8Z#��՛��5B����#p�W�	�c�U�mj�6
f��;�`;��`b���I���~U�nI<���䵫�Ĕ꣜N��{�z?{��[�P-�=X�'s�@�@Z�n����4���\E��?��f�b��Б[�%�%Z��Ð�a)�>v��l5�� IkE!ʑ�/�Vc��I��o�sAu�4L��,t�@5F[6R�T�-O]T�dPB��\�C4X�0{h~�RpݣBXq�F��@�/�8.�l�.%��&~�7�K�D�Q����	
�搘�o��gyP� &� ;��0]��m<k�/WON�X�&�6ܽ��S	���-�p+���S��b�뀫��d�L�k�5\���-���-�,LA zC�,�݄�v�A؆�ݧ��������@Ы��ڣO��nbQ�ad9	�[B��:��!f�%����A�X�VK<�T��z�r�2S+V�0���+�{�Tϕ�O8�E_kLGbs/R� �vG���cW�rT�1IZ�({m�g�^4�E��_i�Ò�ƶ�jz����
���Uղ,��>����Z�=!�8 ��/)�2���`�G �!!�)���oM��
��s��U�V�w��"ذ�B�P!�w��E�Ԟ��E4/K�-6�����4˯)mpܥ�	�<}$bC]i��Loi	�Z�����x�g��꧑T\N�"� �f�'FP-Q�gyZA�����(���ĸ�6�Ѭɥ�����E�^}���:�&�>�<�R���%��������m
�Qt݀%�U�Ah����=��.�8���Ӌ' �yya�Z�{l�,�6��uG/��T$�#��'��b%�d�]f�s�)o��Vw�!Δ���c`1>��re����0R3�8�O� �2����R�8�c�L�]x@�2���,��b���\נ�lC��J��N�ؒt��Ȭ�Hiɖ�(���F��{JK�9�7ye�� �w�Ǣ�k`�V������\�C!W�t=N��Qok���T@
J���Q{9﹌5��t��wL��Q�E�Y
�� r����'����˫���3M�m�Нυ,��A�`*<��6|ǎ��i�~%���V��Z-���K���M�,1��Qf��	Z�<���sW݋�:��4�:�o�i�W�c�u�CF�ѭ8�N��	#$�Z:��,J_�5��nm�t�7F�%�ry[��#`U{$��v�h�4^�	����z��(���Wv�g�$c��D/��d
�<~s�Tm�箒3�?+JMo�0����'"�9�g�c^�v~�wݦ�*BQ���y����T��%�C�
L|�}9�G�[:�
��\"�IܽB��K��+#<�����V�Ԟ��i�o��L�7uKBAw;f�{Ŏ��b��3;�����9�M#�OJ������gK�o���1�4Dr���l�,��nQր�/U�E��2��`St��l�7�?{3�k5��\�jF%�!�d?�Y	�e��6��n�[�E�ah&;
��,D3�NL_D^�⿆j�˘ͦ٦���1�!z��������.���#��0����o�,��f$��ԏ�Ch�2z�L���W�ޱzb+%������Y�Yâ�/��(�X�� h���e�����kqm/��f��vi�����Hf�<�9�j��ZE���t���5jq�s�\�d.��K�g�t� ��֙�<���f�5�@�5��s:&墥���Ƨ���JS�ZZ�x���ƀ�̿��L!�)��誀��e��@l�[
R�>0O�����1��d#�H��Й.��^�;\h�\�����fwq=�Ϯ[�����T�h�\��1}����P�Z��7��,�� ڑ5W�mbN C�)Dc^�v�P��h]�\�O��{yH�7����dU8����Q;^:�e� 0>� ��/;�]D�OGD�>},E��"*�Ĝ��[Ȝ�_��m�<Ɔ�_�Й6J7����'M&�R�8o ����x�������w�=v��kn䘪΀��Q�Ȃ~p�Ak����_tm��Sw}l�Ѓ���W�P���,��['%�.G�W^Ԑ뵭i��
&�:2|�m�l��N0�+t��]�8�
��ߤ��uM�DEJԓ<ey �5HR��V��B1m�1!�i^��R���v5s'�g���*�'�h��Ƅ��e��j��o$\�DŨV-�͒�9�lx�ze�t&��@<�yZ!�8���k��ۮ�i�:��N����BOk�p���i�p��f�rcKG?dj�c�*����M�k����b����m�iQ�I2�ԛ�I�񥇈y�@/�ȣ��zF��J�hZZ�Z|���D��ͻ�5/��/
a������.U�i����8��V���h��nM���B�!���;[�������}�0��+�N��s;�5>�����ߩ0�%yEB�kd;gZ�3.1�0�F��d�:q[�ҷ�8B4OMG���P)��/y�Ԋ�8��|^���tsЫj��	������~Y:���s�bЅO�4YQ�	��~�R�00�zVT�tXlxV64EB    fa00    2970#	Ҵ�j�����L9��Tx�#S�8��lѾY�m��7�ߓ�����bi8cØ�?�r�̑��t����GӘcZ��S������喇旮�t>���'�6�M���	��rZ`g��hW���`u�Xq	j0�X��i�Z�r�q���h��[2�NЉh�K�ی��¹Ǩ��ҫK��I��T�͛A���[�y�x"H�sE6�9�':����(�qK���yk� �R՝q>S`���!:?@��JU���1Vm'$�9[�V�e�Ȓ��cx�9���H-pQ�3II���/�*�90�ҝP��'��������1R �(hͳi���]H��)ru�n'��O�qR !��P��R�fc�����z�bs��Q�
�.�v{����0s�)��
�f� �^�62֏�)	(�q��>��P�K<ُi�A���bK�O������*��!q�U1��m<'��#�8�����"k�j���	󝩵�����N���J�ʐ:q��m�0��DS�O��gk�Z�%���VV{�Q��A�?tʑ4�e�[����M�Gw���IP4�r�=L����
6,L3�01�����K,�fqt?�-|�೓{"��ϑf,�Ҍ�IC��,y����Y�m�`�oA�9B�)˺�"&ROt����~г\"ד���'��c��?�����k���;"ÍZJN1�s|eyB�&���4�4�A���K~U�|���|zQъ8�)����TA�
6�'��@^�d���F]�����p{�~/�p�%:�)�LFq���GRuwQr��������ա������f{��c'1N�q�y���42��3�3���z�sw�	�)���U�5�5w�1��|�1����b�e���L�LO(���5�`�@�Gn��_ �w��U���-8$�B۠R �w��HjmJ諯��Ȧ����tm�7�&n�G��Җ��Ī��8t0���-^�y@��&3t7���6�j�6>M�(6��	>0�؛Ap�,t���#񎙕cmO�1$���9b��@�ϠX�~�.��$W'VcM�m殍'����-��d�_�.��wɥ�d�O>�#�LC�f������/�w9���-�e�$}U��՝�5>�աf��^u�څ�&�V1�W0���,K��%n9oH��G��X��6���eG`V�5D�_��jR�S���أ3�orS�Hr3p>EKԣ��ضW�%�A���=�k�5l�g�R�qSk����� ���ω��j�?��^����X !{���n���������Ho]�"�<����Lǫ�|X.���6�X�c����Ǹ��Z�=���ʱ�eg9��*��㏌�aE��T(s������c#�~��V+�*.��#S�O=�,=�Nśf�Ĥ� $<�U��PT�E��?�I����^&n���vu��<�M�Ә�Q�RR	&�bٲE�"L|�5< ����� �p���>�v;4���C��2m�5WG��!ģs>�[k13i��$��/Pb�жV,l<=�#oS��1�g�|kH�i�h�?2��0=xy��U�6��^�єYƚ6�k�ג$B��"�iqA��J=�H�x��ސ�.m�R��D�_g4I�JKAn�UB��?�s�)/�J�{ ��z�c�5�A���,S���VXw>�Es|Mcc!�%6�]�4�-G�T,T8$!��0����|�[��v�fj3��=7c���#���gP%�3���y6Q�
�1� Vr�8�:d�ž�������1��}����n��4-�৺��ʗ�2D6����DgZ��#�I����*6ƲI�N�n��mz��^`�(v���)J�y��S$�=��2����|I�3��k:���Y0�x��b��r��H}�X�P����\Ar>�eCo�.���lU����X<�rq%k���Aa}p�Ee���+8��'9[���$:���ҌS�ϱ������}4]�b��Y��mB��,�m�j�=hc5��o��F^ďQ5^��]A�H���i���U�	a؅7�&�$¸&ٓi=|�ɟTL�Ø� w��K�i_1a���Q���2Jr��b��J�;�,��N�y�6�!��R>y��[���� m�[�N 0�?IX'�k�A8��.��C;�N@)E��L����b�+�pq�O�����<,�a����*�\Zs�ƴ��[Q�����o��!�b��ǲzQ�ߌ�&U����]=9j�]hBd���H�j���s�a���Z�P��CX���q�<1y6@�13�w�V�g����z5S�hBo�I�ݢY��fRp�䂰�G
@���R���<���q���2�04-��R��ୟgi����b k	K�q���Gx�:�ыг
�̦�J�ܢ��6�+Z��As�d��4�ru�c>��u�&�[N�/��� !�
O/&f÷�h��nդ5 O9L��K�D���
Y�1~���*r��"�?n0����ޒ6��ȁ�\Ԍ�ju#Vu:���:���]B��/??l��c��,���[������*�!$K��� ���.*%�<���*�j1o�ō5a%K����X]��e�b���UT,D]��:�A�{S�~ �[R�U��J�.&7�5��tdUt�9+��޹���6�{�/���a=bj�@��Օ ��z���*�b�W��^Ar�$"�J!_��������9���^���j!bMށo�l����a�?{��G�7#��]@9y����R~��+��Ad�:�d�6�����F��^���E�����$��_���om�2[7^)g���Z�Tޜm��n�hLKvbnHd�������ѿXR#�N#4��I ���	��w�0�\���3u�!�F��L �X��o&�'�
Ç(.��vw��*�l�*h%���b}�v���ޤ��FS�Z�kk�9g;����{���9��0��h�㻛��7`��|U�L]�B�'�������l���j���gN���}�Yr��%�i�_�9 ގ0ÿJ�}&��O�`V���-�>����`�G�M�ނ=�ɢ~JDVo�?��+��(�%���)4˱s����X��'����A=���eZy�'S��$��9��|u�H3;R9֓z�����c�٥8H5u�f�-�I|����KIq^����hkq� ߰�c7�=d
z�8a���}�����9Rl��rB�e�,f܇�h���cS1��.6mG-+Ӵ�!;�(^ws��?��'��|���e��2Ng���������hl���')eV�-m���Uo�n�jY�JJ��/x��KO�:;�Z�wik�B�ֽ����´���l�8�+��t@��`Pǝ9ɚDp�z��,)�ؙL/��� JЃ�<1�\e��.�3^_�pa�Q�I]�� �� �T>z
"΁i2]Jse����Zy�L��C�E��뇆�]��>(��Ը/׽�Z�NǄӳA=�(��Z*�2Q�"�C��0�����5\Ö��#˨\�w�����E稽;'<��\n&O��䒟'n���]�x��]�Dy#��h�J�b��Xb��'����N�[�s.m3z�3�Cv�k�N�Wc�r���I���UM#�|�F����H�� 53�$��֙GU`�e2��>9�w�m�I��Dܭ����X�Q>o�z&�@��9����#*�G>կ���UHE���t�^���󫮭:]M"K��@���0�*Zӡ�~�)�!�,�*�k�?s�S��. F8o��o��,�XφsD�a�E��q���~�|Y��W*�B-�h5zk���ٮ���Y���s�����w<#�4Oc��@h��ڏ������k^�2�J\�߻�J??cߒ��o=����s�9J�99rB���䤟�L���l�o֭�}X���-�`+r�<oEc�o|��>k�1���}��%��o7��s����YSͿ���� ����J&����S'=��9̹>2��2�m�e�/��{"�]��*���L��]a]����6:�^kef�|`��Y;ޯg-�6(Ј�\��n�Gw.wل.������}�������l_��K����.���(�̖�;&~ �(��/?��d/9����\u����F�r�h��6��3\Ҕ�G���FiFT���Ӟ���fAn���W0E(3��=�j�>�@�w�Q=#U>k���I����P`F���$��#��}���@�u��+���UN�~h�/I�Z�#��`��V�����1� \� $I�_G�9���a^H�^�p���#��KG:@em��.s����e�>�%-���	>�lm]f+!���!kmo^�~	�q�7T=݌M�A`*d��z@� ��[��������$�&"ħ�����k?��nu�8�RWF��TD��e������F�&vL���&���u{���>蘿W@_�&���E����uL��|#�f�$ܟ��'v&�w�Y�X�!,QJ��� �]0Όr�O�>V"N#~�j�
(dO�{34�t��O�JV�����Q�~k����	��])q�H��MIڜtN-.����c�}�vz���H�?�\3�)�;�h�n?Fq|,N��f��@d�#"�6������5D�."����V�l�uL��j PN�����=�51"�XD��l;�j���?��W^�Q��P%���G{Y�����L�z�M^߇_��w �'�b�qI����끺�$����8�u�%G�h��hB���~�F�L,bS*E+������>ى�R�K��R8�]��/�����|�����-+���9',ŽyR}�+�I���`�CLA�J����`>�����_`��ڒgk�"X�a{�x�&�9r2���::�S�/�&��KE�c{��Ry��������N&ٝ�uXQ8�۷�ʟCl1U����a0�
�W�C^X
wIP���YV��ѝ���,KI���#5�U&M�&�_��`����䗬Vf
���%��	�W;����ET��`(w������(C˰��a ��kn���{�R޵��ڵt�t���%2�~Q���P�e��n��/���K��Ɔjx���d x
-؊��n�V���#����>�sv�!e��uU_jj�0�e����؜�� �N:�6�s:����:�O�;,�(�!���NT-�9J�hk3��xa�a�+�ץ~�eR����陡N=My�����@z>��rh;V����h�r$f�����x)i9���G���l�ɔ�b���(�QQ� ��тO���bL3_����%)߁'���x���Y��xU�����7��iĖ�t�{h��T���Q7�} P1�p$_Qv㜌�W�Zģ_w���b�9[��K�˵�7�k���vWh4�)&/+�l���nԯ�8&/��Mx�Zx�=�V�eR�꿉�s��F������{�O��T���Rj"��kf��.k]�-�I�f����}}���iږ4m��0ҘN�j��-A��ܩ�,�S�J`И�NT����#�b�ΰzLLcŧ�-S��V:1�l:�ɡ��Q4�"�j��jF�4K���\ի�N��X3r���y���왰�6Yn*^L4dX�S�����׀�8���j8���p��d'��D�ś���=7�-g,�>-nu����2��'������G53"�@�:4�O~g��bқ@�C=>D4Q�C����?�+���Dl��*pG��6�a~��_��
7��,�}z�K+z���=7Cj�ŉղ�}�Cb`��t���k}}�L��{�r]:/���NW&EVO�y���0Tk�p9�d��Q�9:��q���^%�e�&l
qѰ9�ʜ���R�X�U)�¤��/,ݘR��fQtRh
ɛ�ƴe�Wt:U7Ӕ]Bo.�jX4$�~q� ��AJ?=�����QJ3�;���H^�y������-j�Q]�<|���	�B��D9�5��DK9��;���G,�����X� -;���G>���\��Gxq�+�AE ��s.O�F��x�\�X3c��-|���K���C	/�U�\��_G*� �(�ӭw�����l�g�QC�w	���@FD*��YqO���Ȅ%�]�R{ �]�K��iCq3�v|�u�R�,\%�������S�t5����E�2��9u���w ��Gxdb�@gۢ#�.�⹝"�"fB]�E哑;�g�]�A�4����Cda%�CU����Я��mk;�S�����ʛ���"I6�bס���V%x_ P�3�=S����4�>�x��l� �ǅ{��t�7���V$;#t��K��J�Y�q��*�]f§a���L����$!�na�Ch�;1�ӰWYDV� J����ιI��l`a�K	�d��ܫ8/졅+l������-�1[�ī�����Q�~�SI��c;ɐ�ޘ���b>iT��ӂ��&"~�� ���'�x[�_wt�B�EE�[]��l<��dH�oZ[4��oo�7����A�ʈѧ:y�'p���0�B����lWH�?F+F�6W,_ܵE����?��ro-!_�s�
6��"#$�ȾR��/�.�4�&��5��r��Hi��r?֏�Zߴ9��@�p���j�$��uQ��u���r��� �ݧ➟Z�ȥ>�#����эU1�=��K�����Y~�O���@��s����,�W�T�������y7=S��|)�&��zg�\�i>6[O	�f�WS8�Z��}L-�1#e#��c"q�r�Xa��?�����00�+H�Z	�	N�+a�W��a�(�`G�+�qj>�ڀ'TM9�����cYKY�C�I$J����_���0g�FJMuĄ =����g&�5��:�,�h�t�枧X��\������w�b#�[�B��?+��]�Ǆ��&K^��JMl���U&g�@��ǡ���!p�!(,\2u�����e�������4֝\PdT���6�B���m{��?�5���3e-��A���4q��;�ؾ,|쇽�L�%E��N�$T�"3zbl��3 4�(C�0B'yȂ^Y��*�l���{I�k����xh������a��ܧ6n�B������s�EXP�l��-<tp_�k�φN��� ���#uE��u���=K3�!e�j{��k����Z�qH)ZhaMa��5�/���@�ZH�Xˌ�Fi��="�T(�
ò��������o�U
����ؖBl�.N꾦`s�F���$�<�h��g�9��nJ�i,�?�s���˽���/ʝ�����ۂ��%q)k�E[�i�Hn���"��~��Zl �`?�3v�㶍�����d}�0�؜�_'�g����sgU�GTP:���s �����[P,,����n����Y��Z��}%�����EF2bE;	�K��&+�ghR������&��`:q��: z)���첶4�t�?�:�G)nf��Δ�mB���ύ��$��<�q�'ҝWN� �&E	����p�Cֳ.��h�/b�a)�;{Лi�fahVG�aj
G4�#�Wv�������C3/7~�N/e�H�ݨS��[,�9�#����1Y��T����\�����\A�(���4�d��{�8X�0[bs�o�O��1�D�_�\��z��9]�N�*�[�Mz��ܤ�tW&��m��1�^�#W��l����!�l��5�ב�e^<ǖQL\�"��m�����vy��Ä��/�s�D�)�/ֻ�f�ݽ�d/�����٢{n������ߙiԌ��gB��4�=U/�P��+0�1!:�����6���Fk��14��>�M~=����_���%�����8�).O@�ֿmY���!��	78�!3�����p�͍+?��������n3#!�}�d�L-�b�ǄG�ל�}�}o�mE|��XBV�qGPqb��:�@��˽�s_�R<�f����Ef�����J2�M2�\x���J�e�<�~D@�
���џu(W�n�y?0Q�7�VZ��yL�Q��V`���a6�����zѢ%����%�Mw,5T	U^1~h���#�H����Κߝ���l��-A����\w,o{�Q��s�-C@�n��hbpA}�i$������l7�]&cc��j���E<���&RLku� RV�i٪�EEB�:-�I9�-��&춎O�"�/3�B\Q!o���f���w�f����@��e�p^Uy��
�p۸�K�ך�odXp�ܽ.�3�M�NSo,`�9>��F;��~��a�V��7O[L�6\ܥ	;����a	S�b�L}���7'.�Ow��˿r���ISe��Y������l��O��%���f$�A�%˘�AU��A*5E�B�t�o�f�u!]z��Jb�5p���)sk��2a�	����G�J�R�޴�]��bud������o~��O�`���2I��`�l���C�P���t�if{K�k?����#����S��n�&�f$��"Coά?��K���`��ӯ[� ��lm��Bv���\�]wїXM��C���b�aJ 2�1p���tww�l��0H�3��&��8Ʈn�s�`��(�f^�Z�BZ�0��!�
�6$/��HTb���`"�D��M�$���dWJ�3����l r'G�����L��5�uw�gY1�xƙ��n��p��4>L)��XߣȦ�y�1n����+n��9�h���aK�����wcg]�Ȅ�"��t�����S�/қ���R=��ӑH�zy�ie���N}ab���n��ܓ�����v�'Z�y�z�������y����E��yv�=Kݎq�,� 3�G��PB��8Ov=�s����;h�����*�MT;�$�?��Zo�əaI�z<S��8�~�|2j�_ל����ⶓ�B�+9
&��}�B�_�s���!b ��_���<���nlP,��z�UuW�aOP'�ѕ��z�6˧��;Pv*�#�^~>�ﶡ�F!��\��֭��Č����v76|izLR���i	r:`�$sp˛z�3e��8�v��ͥQ?�ɓ�!Kd4g���1���cl����g��� �^���2�A�p�;kZ/��m��_W��1�K����KL�6���Ou���p����0��e��n�jέ�pV������R;<�N���������4Y��#U!�v��s��F;�#��>�I�ʘ�B�x#�20J!�� �L]w���i<�#I_�����j_�E�˚1zdS4p����[����\���*Tҙ��O~(t�Ca�sM8%�lXKA^�I�N�t�(����Q��FȝJ���h����hр�rP����0��-t3<�0@�G�bT��Pp<�/�T��)�o�3�)�|����>]E�p�z�ꅱ~L�����0�$�v�U0˹��`���^n[�����̞s�s�Y�ռ��[mr7�C9��VV*�ه�z(��*>ܠ[��6�Ы�i�	,���$�e�1�_��l�TL9��y�c��đAfg8��zl��x�<.�`�Һz��s-߉i���o]i"eЌ��Y�����^��UBU�w�N�0ux,>G�'���A"���V��l�2�W{P�[�Lrw�x±� ��s���@\��V(O�V�~�l-�	�3�2�ڧ�dm}��1ɢ�Y��X9������B�8�U����p��OJlc���Jwӗ��v>{?�E�/�E�4��*(F��7ӗ8�|+���/J\�u_R�h�(��S&����B�0���z����[+;�}̢�p5Ln�4���%��%�v���)�(�aFS�;֪D"�vV|�&C�vg��n�T��Ĝ���i��^Ø���CD���V1��������'�\���A��O�����G�#hىF�C��3q�;P��΂~1K���� ���V�ʝ�;I��Q)� &�Y����<%A�,?�#���$�\��P}�B-z��/�J���4u(E�[��R��$���Gق�٭������fs�r��"�=�T���lX?��j
z_͙M|!�v1�ڧ�Գ��n����ːR��v��a��p�f�l�Vo�8dv�c�T�A᭯�>y|����R%�%=D�⟝I�F��Bq'}v(����Hs$9s�
íl�U�<����[7_m��+@�Wģ�8`��	�M����S��i��!V�|>9�%��V�R��(|����w�}O��y�%3�T���Ed�`��)��IEyf�f����P3(%�����y�;	��\>bUf}�f�4"��d�b��zb����UEI>2<��ь�*��fu
5���C�A���ynGO]&�F���K`߽�|CɅ���l�\�`
/f��Q��jU��j��/�U�����TY��c���>_|>[��O�\��`*e�o���� ٍ�m%_.2t��&B�H��۷^��O�LXlxV64EB    fa00    2a80�rK� � 3�����qa�j��i��$���x����%��O���R`)U�X�W���bD�=/����hZI��/�����d���@ւ�ޔ�)&����m:�&V(<�!J��Cp���d����O.q�5��W�6Ϲ%9����+{��#�_GvCF���Ў0�]����w�mp�-�U����R�0	؀/w�����2�q�� ߹5��@7��H)��s����L����N7�?�k�]+�:�:f��YNUq��̘�eN�~����'���1uiM��j2�>�^H�p��8�S*��O��^)yS@�^�C�@.���N�>��7��	�pl����g�3��Cn�>NgHl`{�5A?:u�7�!�����z�K����8�jf�����u��4�Q���|���+�	�- �� 8�F ��� S-U�q����R�^�$ߌfa���f#�mZ+���!0E�E��e���#ȋ���Y�)��d���)zC� |r��Eh��[@9�ԥ���k|m�.���z [�طQo��qS��d�l�~��~�����Uoo�a�.V����JnG�hn|�e���Nv���1��v[�{�����3�ںb��B�@tm|\�!Թ�-�s�j�T��2�&�O>f��y��#lgI io�U(\f��	7=��%y�� P�åN��{��D� A�VŤ:��A�4�D��߭5JU��$�,�b���R�ϭ �v�6r!
֩~pŨ��X�'Ҩ��T��0b{�K��L���ʍF��lv�j��w<��Z���I����6
\J�gu�=G�]"�"��t��袰�
(]�HXg�W���Vnr�Ox�Ҭ7j��94GzM���Wѿ<�b�@z� /�SdTL�Y>���1)f�j��� ЍZo�虐ɮ��yk��P��I�ȝIQ���=T����.�/,��G�����D@wkO��7��GV���v�_h�R\$`���U=+9�A/�����1i޽uM7q2j~X�ȞY #�����F�}M朗;p�B��_��V�⸫4�2��Y���r���ہh<q�c^;J�zܤ���a9E�d7�H٬N1z̄^d�|������J�=�_h�]�����	7KSq��M�w4|���s.�aa�s�u<�ݛ*�Db+o���9�C-6\�����jk�&�y�V���td�N-��[����GRH�-M`��ʚ?�a�8�����J "3a�3K�=���ng�CB_ǘMG �5�?f3X�GФ�H9�}��2�K��/]y��=���e�H����D�YB_��=���D����ySL����^0]�wT-9�(�ESEN�.~Kl)�'@n��-^E����J�VtI�'��`��l��@���x�]�.�@�w���Vf������W3\�
r�b$�+�̓!��TWlvZI�DV3���eݷ�1!�rGł���P1�Jy�>oL);�6A��#�g�9|�����6�>Q����>)!�3���]��҇-�������ǜ��Mr����ae��S^�?��)�GB�^�+��� �">��b�y?Ϲb���@�ߢ�(px�O��h,H�b?�:�	��O�q��m���S�fҍQ("C�z�},Z�ܤ�����f5I��,(�/?���90"Fs�ƱU��ExW|�t�iZO*4_�u���o�d�(�����@*�+��9�p
:�����B���Z4�`l��]��@m��Qˑ��`¾&��T�u�$8hB�$77���Ca$���d'(wypc�2�4�	Kv+� ���D�z��G��hn���-4�gj(1�JK��)W��Z�ك��C&���f��`�˸e����&���3b��o��;�t�Xd�~E��Ѣ|#v�
��ĢƉ��ຮx{S�C<q��H}�n��7�z�JJ̩Ԯ������P�������D���5T/��aJ���a��r��:k%S�pZr����e�,+��
r��$�˺y&�=8���:%ǌ�n��wpu,l:}��a!-xt�}��h�se�ϕ}+�k��2�?u@���{wW������A�dU��p�0�mi	�V��ּ�({��&����7v��-f0��1bp:��h�mh�	g��3���lU$��k����+X��!��=�'�GϘp�<d��3 �#~<��ق��FXM �ă�J�B�\la�&%��:�������~ǒ���킏eu�����ҥ�l*���dK�uuH'NS�ɱc�ҿqn[�vy��xS����uQ��˜&�h�n;b��,���0r1z:v�i[��L�,b3��Ƈ]ځ���uFH�� ����8�*O�6��nv����͵�W<��Ι+J�FԔO���V��2�q�e��?���|7ש�P�aodBZk�������g'lc/#)��ԳT�l���V �'�de�W5����#i��k��wп����NБ3��y
`�/N~C�����[@����|���C!f�F���FH��z��75&Z�z'����)K%� ;P,�� �4��Q�x����=^b �=����pQ�=��}�P�ۮ�e;�5�z��)�f���������/�>����,gX�.�$��a$'�������)#W29�3���O���	/Z�vi�n�2��1�7�U.�ۮ��<���0���Æ@��n"Ri����4\�p���,�#�rq��i�Y�;V�_}��dW����[��)��54����4Qp�I7��]V�+��W�v\�oa��`�-�f�7��PU83���� 0v��J��c�=�8L��8���@�3�����!�K���摄/�Y��t��s*G���� lU�^]W�I�8�y��0��uvn:Lx˲�y@�.N�^"
}�ٳ���������	zn:i���5<�au	��^�wٟ)7��~~l2��#��lx1�a��٧r��(�n����<�������Y3D���(#��u����l��,p. �f����N�,�a�.�3<z���c!�綇�_�����`�5؜Qm���86�F�{!�FM��k&��	�?(�(��ަ#~Ğc���X��x��8m���gH���_	�/�GC��˩<� t\�AU����L��`aP�@8���zԴ��F�Ъ�l�g3��&L�`�f���Q�;�<�$u~�9�ǝ�eru�5{@�்�Q���a4Dk2Ng��c��A�^�)nB�'l�:�38?ь�PR�e�h��Pj���"��0� �͏�b�[��,f��D�a�K�HB7��!)�O�LX���x,^�y��F#\{U��i�B��H̪�9P���oOĢa���/7�PY�t$�U�4F�Lś]A��Df�s�	_-)9C�qA�+a(��I֢�?1@�	��Uƹc�&��I��3�<bM�z�ǃ�8C���7d�..kc�׍Za���E͡wѶh�Z?���C��[;��Ɇ��Oy�-����#���a]�<��̢W�����ϼ@�Q��C�.3ҕ}���j�\t���/���˔\1F/R��yhM9�BG�Ӫ,"��������Qz`��=B�[��*_���֤��g��t?m�?.H�3��|H�a�wi	�*�ɞ�� N��QE��$ħ/8k�V�q���� ��Q��a?m�iL�N �н'R�*u2���q8����3LFbN�+W������UcK :�lPֵ#1�@�Bl�$�d�\���/�v��+�&�����Y����oL�����IY5L�G�n��r�eY�9"��oE�I|3�~�<���Kn�	����Cղ���$?U�y�`)�y��9����7�mpL����bm:����ݒGv����\�7�_���6�Ҕy����św����"�+>K�魚aX��q�q��G� ����/�t7 ���ǆM�k�=s}�C+���JWq �3�j�^����PL�k 1�h"�<>m���
A��;3s.̹us��?|�K�]�щ�>'Y0y[���9�i�y�od�po�u���\����A�6kA�O,2�/0d_
{��$���Y�)��{T,+�-H��ț��v^�؆y��I2�rmw�u�(bz0=gk��S�M������{s��/�qa��S=���yy� A[0�>�'n�!�j��O+��hS,�^���M��[�su�X��m��e�m�0�A���^�(1���%�y;�hZ@��|(�d�T4^�qq��~�M�S<p�Km���BU���ef,�qs�4m=�Ö~��Uy��f���
�)��w�,M�&Rhx����O�I�Xx� T��* �NÆ��7��/!�'�=D����l_��<%��ִ��3$�G�]"���<�uLEZɍ�L��`��4����x��p"Si}r�ǡ��Ƭ��b�>����`��s{�SyeK�s�m"6���azF��$>h�Q�4��6��B޴7o�wɹߣ�q���L?x$����D�?R����ơ݂�����6��t
�PC�½�(��i�=M���@ɀJ�Bv����1[Aۂ�)V��P�����n�A������N!G�fS6��s�t.�T	9�tSU���:N肙��$���+�ܱ��J�fOƀ���������b�~��l�>v��/�� �}�
F*&\N�tƐ�WI�h��ݺ�Ԧ�@@n*���#��L�^��Ec�'�T.�d�"��s\	���% ��R�0q�&����������~��G�Y�8��^y��H8���Qc�����������J�{[ �?_M���e��j���~ء�w�ǽ�����H6��e��L�QJ��`rIcM��6{�l�x�s���P��P�n%�z-�H%��ۂ��~�쥊SBo3�}A��E��tF�O�����we�^���@�ma�W0'���칽�VD	n��1�_(��$QxF4���|�"�d�U30�Ûg�s-�޲<<X�`yi+�腫a���j��A�!B���1���7�x�C&;�x�\!AeuoAI�{����][�,m��q����!��y֟��5���
�f�?��E�6MX8ʹ��9w�o]���w��_<���!��P����7�"�)j�G�&߮�CK��z�~ܶ$v?E%�P�|�kf}��Fa*<��*�
�T�Nk\����M��2��J�^�_��'Q�}�]���;g!���Un�+sp�zKZ�gG�������"�vp����zݡw|�j�}e)i<�
�z*S��mJ�ٖ�*�@Y��@��~�"�?l�jT"�������v��?&,�MKq /:��#R�<ڗ�П��esq�����i�`�S����)&�TMDn32�M�b�n#� �N�5w��8b�����E�ymy�4�0��6sRW	�mG~i_կі��)M�g��e��P�ƒK�Lݗ�б�a���곢���g(h}T�/ǳ>�����.��Ó\� ��?lA2r�?�Ζ���
�=����(��×��:�~0i�{J<fp�Ќ���q��s�0�"��tۢ:)�M�w!?n�#ck���mS��o��U~S��& �Έ�4X�w�//jҲ3B�	g�%�DD-~z�@����l"��ѕ��|j\Lކ��ϲ�$��f�D��S%<�\��ɢ�Gd���]�V[�c�W��Ck�t�`�('��/���Dy��x�	�Dvj9��]���}��k��5��p�.�+�,4��7c���Y�R�?�ኺ3��I�%[�nR:�1'��jS4�/�,wr�S:[FPşn�գ`XisYm:
:6��)鎞�e�IH	�ʞ�\`c��������3���ǣ���������B}�����c�*D��`��d���o�MwI�p�#a��=v�<�p�45��]kI�c���r��Ff`�h%�8D����l}��)����NC%0���~�C��G�/�^F���W5N��U��Qk-�މ�x�݁J�HFC�,���^5�K"^5	7�.�r*Ψ�^�v$�O�u�_ B��a*ʒ����9�AF����T�@�����e���'ض0H��I�~7EM� �LHs��S�i�����{�QЛ�0��ߘNUiI�9�
:9@�ļ����4��
%�6ȃ�[��/~O��;�����xeV�+��P ���#I1|k{�{��h�d3uR8�w@!��_jǐ֍�,��>=���i�Kqr �gn�ל-ܸq%m���3���v�6T�O���|�"�O&�o����fz�T4�����4l��=���l�db�����Q�j�i�2wB����G�3��X��\p�`d!1���q��w��PnaiF7���Cb��4rg"Z_�3_>�j��e���n@����33��rykQ5(.�5�E�W���G��ޖ;vt�_��k��Z�o��C�j.���4�� �C�U@afak�1c��d���^(�͢.Z�F�������g��Fx�[H�~Qh	iB߽v-/��[�����]Y��Ȳv�$٠�kV=�k���v1�bUFg᷼�������)��"׾��Lp��_҆��@,�SW��m�N�d���h�*�����sfJ\|����/�`⨴]Q�y' \������w��E�0�����貥)xl;��`l�J���WViB��f����<wpJ�1�9�y#r��#R#7X�-� ����ɍs@^� �CSu�s$�IJ���y����S��Y*���k&�����`a�6����7���ї1���+��&t�S�ի��m�&L^fSS-��ԯc_ќ˚��<��ZǡTP��I:=*X�s����6 F=C8�ڹ�����jcF��D�J#��'}������X ±{��ȥ9�ϓ�~׫��q��"lw]��w@�S�����N+�W������6.Z��+oX}`|��ۡnM��11r�]��Q;d�����툭֊���(
�����ʁ�>Pa ��n
4����W��C�p3���'ڥ�C�2�󭈃 w~-�Dա1�x��@�L{*(Hݯ�o���]��*8�g��Y��H���H�}�����>�?eI0�����sR�U{Z���%ƴ��*�7>������*¹s���P�?��T 1,���vb8��E�S���[���̡:7h�^�L��d��(��~\�Wt�ϫ%�JLB���A�"23�K̵��S�`��\az�F�S��X�����F{}W]��o��%n)eA��o|�W�i����ew5�{VL��k�省@rz:�\���`�����3���J�?��:����H91���┏���G�
ɽ=f{6 /@q�`b!Үuw�2?6����d&d �r�l��~���p��󡋢�U�s�,S��/�:��=lw�a�5������/ a�M���  *1�4fyx�]nh�W�!���z���@u�]�����DS�2~8i��X���~�+w�gf���zy��b����4o$���Y�_-����ۯ4_�~ɵ�3��HծZ<6���yC�L*<�Z!� w���*]u������ٺ�;�Cl��]۫ "��!��t�畤�U�X�{����ޙ�
t~�hۺ)��c����G���D�q�թ�uMʱ�E�'��-2��~ϔ�!���"��v1�j�a݋%�
5|��-I{A����/F;�=�TF�7	⊷�g�,J��YvR���n:�pec�}\)YmH��{�0������ ���*�R�a�lR��������@�OZ[���k�� A�v,�����]���ܘ���T�byR��wn,��!l��s�1��݅rt&̅�"%w������f����5��)��o�� h �_����C*�F�鈦*ͯa���^%_��TRC�R-������@��R����*�PMn�t�4t���1VO3�������=z=�����Xû������\֋;�H�τݷYlpDA���l:��XC��n�������A�TM��JR*����j ����^ŕlKc�����"�EcG/�L�ɽTeҤ�v0����c�u�=�����	���:>�
�>�	�r*�j?*İd��&�z��Q�[f%r�Y珄.aK���O����I�W��NmjZ�u����9^���]���d��2G����!��G^�F��gp 1�y.��R:���qM`&qFq˓�6LxE�ޙB�1v'�@<7x��{�!��m$���s���Uo�z��F����[�%ۿ�o�,�u��LG��:J��l��7"82i9LZ� �}OY����գ]G�Y�hˌwi>�h��ͳ�%���c��yf�p�b�����Հ��q�I?��9�z�a����hK�\�6�̎�y&I��n�4���Ԣ���/S�W��
��@:=�#p�'p�s��{����т�[������&���I��=��e�����r-'���8k35�4E�����&��s���6��	;x?p�n�D���Q�&, %eg�ca����&*�}�C+���6/-��{Ȗa��3��B<9�/�-�'�Cu��j�O98���i��>Լ/����b�vsv�3�al�∍Uv�2_�eYUl"�JH�Z���2WO�ׁQ�7I\q��K��:#�w=�4��Vd�zM�#���Jw�R-ˍ��;�ƾ�LQ��^�^�"p\�5#�� ˠg�j���z+��rԽ3�;ӭ�㸪Z�y
M,D26W���z�>�%�2<=R����y�"������o��YQ��yP���o�n�z)����K�#y�9U�H��B�0�, +1��;ڥ��LLJ3�b��L̦�$�oX)/���κ�F����f4i�C�a�f��/a�(�߼%5�!$���(�Ʈ�rA���F�b��t���+�N  !Jxބ�hຎI��+L�6T�U^ri�Bbb����G���t���u��>OT����}��������]�h_�*���'���v��/�/mh�bK�+���Qa���w�S~���n ��!7#���w� �وa�zp@��3���W����1�g,��6l;�CN�"�\
lRa�e5�JL��J>��`��T�s~�2
<�?��0�M��v/]S��Lm����ʬ�n;��IJKs�S~�����Sjz�g� ��k�j�ǅj�9V���AB�s�e(����5u�1\������cT+��Kv�o�tm�HE�t=a�R�k!)ƥ �WO��c,���<I�=��UIP��s'�Q��-)�X��+�ldo� �Y1�2Ɨ����2Y(H�G��H�Uq@L˺-,A������[�:?�tg�������G�(4J��|��MfI��j���(���g0�l�me���Nl̒�Ќ��|1)ҕ�����X�.g*�u�2������f��gqM��Y�}B�d���KV��p庀��|�2����6�{�S�U�_J����=YG��WB����3=#[h4�y��þ6mU4E�W���<x!��L��N+:Y�?�Ƥ,
��=O�i���ʙ[0j�䳟����$�ّ�qV�U�G]�_Mnȷ�6�����������d����Hř�]w5�A���-�I���rsЂ����Q��s�H��z[��3�OE㥆�6�Ҫ�V%�;����]DY��8~6:L�oA6q��%��b�����,/sd�"�Z&"��<�*��*>ͧ�'������o�E(�S1�]���2×���'}�����AF�����0Ti�wc��_S:�]���j!%a��k�6���z�Y�|=I󥏍�r�'���_|�.bT�Z�Q,��W��.�HB����"?.�Z[;�V�R{9�Ľ���e���T"�@g�
k���ڋ��#�2Ʋ��o���׎Z��`_�:nt��4��^�&�n{��
yf�{�X�7-  e۰G7���ځ�g!��P�9�Р�ff���ə���GZ���]`�����%�����2=��VĂ�����h=ݹ��rN6���(�_�y���'��{�'D��3�7M�ӓw�#�n�<D�o�!$I����ĺ��˟�9������3c>n:|�϶��P���o478���h���(�<_�s�#"G�Ϭ��>ט�d������w�z�B���G�?�=�.�ߝsv�[��|�����8\�6�`�| {���t��cv��}�	2i�����:�<.�fOK6z(hnØ*!�¼�k2��U|��\ZP��B���{A#$�RhE�&4���F0q��)0#M&(�x�v0 �B�I�- a�B�#�7���L�Пd?�d�ʧRdx �Ay&l,��%���*�.-e<ߛ����"�t&+�/@㻆�=�Aŷ�6`��%�N��='�/�i�^4@�����j��,��'& đ�KI��k��-h��j� 2L��L�[��"��̱�c-��G��c���T�(��O6DRO��ӻ~�0A�Sf/���?�L�5R�;�� ��F���ȵ�D/1>�xC�/��v�ٟ�D�8�5�ڪ�K�;��F�Ll�( �D��pr�F쮂�g��a���3�e�������x��3hA��9��$_a�0�Z�M"^XlxV64EB    1549     530r��>\�E:oh�|J�/8pQ�<�9w�X%߹S��{��7�Q'2��ӟlE&�^(D�]3ik&�y��gLPj�i������3e�7p�c���:�x��yↇ'Kز��dݚ@ɇ����w3�y�;7�ƌNFaHϓ�c�	)�~��Xi��w�M~D���13���瀞��4-�.l��:	�c�.�U��0�0dr�E�J7�>_D{c�|p�=���K쉹�tX��� @u�	r�(ð2Xh�9(Iuue����Qk�t>�Q,��C�G���$d��e0�*Ӝ�Avp�6<��X��$E��5y���DP�t��\��
�_aЛ���p0w��������z�:�ޡֲ��N�:��>ժٳك�׷���pD��\��Eú��]��^}�'a�}�he�9h5)`�u���C�%�����
<��<�1�J^�JjTOpyt�q�I��BL�s�d��%0n�
7���1��5�����������i��WJ0�g2A��D��*�(ɑ
!����jr"]C�"�&���O�Ma�����0��2�����T)O*�2眹����Jn�gZ��r�����q�Q��`��j�9�Q�B�5�ؿ�6=�CŎEڹ��`�2�/R��d�~5ƊnN�6�-�t�����{��5�x��I�s����S9��	�)�5���S�V*v��$c5����u�r�w��ִ�9�pO=��rdͥ{0�X��(ҫ7�=̀�ǭ�]�\�X��|�=�/��r#vg׹mT�u�h�Ǳ���~��R*Oi�k�}�=�2�'�	;ق�~�u&����h�JH�;d�#���d��y|��t\�2-��wm��q��b������n��*�� gb f0��¢lLi��H��<k?wt3��;ϙ+��t\���҉}��dc�C{%W��p�l6�ł�
���p�N��b��#X��}B�8R%�mF�q��KV/���Ψ��5�/�{n��ѯ��Z��h�Ҹ?�-tꗫ>�a�KUJ�o?	2j�qFQ�����_?� jNr|�y�͠�2��� �����x�;�e47]��*a����Γ����?�_}wUR)��#�KPk��������8`��`K�N��6�؜����a��k*pmb �q��b�S��8%�p�eXo�_��.ޘ!M�eсZ.7�Q!�����na�j�YKb�C4z�ms�g�ObD�>�����<=��������X�yE#�a�#7=��dA���v�#_�;^q�#��~?�2p��S��	8�A��)'�"�Z>��e��`�C:���I�6l�nbʿ�;�(#u�v�Q���J�,TL