XlxV64EB    2232     ae0����$h�9�u��/����s:���->�/�7*�}�"Ryw{��~H9�ii"�?��$XF�38�X�A�2�e��V�Ra��!�m(�/|^C�w�[1���6�2���ѫpv��M��� ��_�nQU	ؐ���9r�]�o���a�-%Y��yZĻE]����S4���XS����'��1v=BU��
O����jW���n��?�6k���q~�:\#T�)�ƌ��q�Db��&)�>�@�c����;�(W׵}Oؖ�� P��-�4{4������?����8����{;��Ɇ1Y�}\��⊧��8�&S�gÍfJ����H-D���Һ�]Y��oq$,	�����;��C������H��5��	M���2�ڐΩ'�A���i��R摎MM��"�Էb!ɢ��t�󢎖,#�9ۘG-=%�k�mK���^=A�#�#�����^`Ƿ�k0*}96��?p�g	�IN��e͘��@�7�nN2׳_W�Ģ7=4���EK�ȸ��8+G��M��{?�UkD2��jTC��6͵�9$;��`�g�
��	�;�A&]�)�� ���' �Z����� �F57\�>��nb�9��_Lۀ�����㬺�P��%��y�1�p�=��^Ybh��촅O'�pB�qڇ�ώe���o�Lo�������mq�BMn\%��X�u1��o��2y�����X����!�n���<�ڟd���@m��l�pQ
[�6Gh��=�*��"r|�d�fD��	��K]GԄ,J�'I"�3��M�8w�|vib�����Ha�~0��+��5�*�'A�-Ů����ٯ�{w{�E�jX����Bn�s��� Q�xT*I�=z*�c�Zhch��E4T�;��_d䢱�R^�x2'},�#�^
��DM���g}˟-c7Й���Msc�;�$���R��!\��}�C�sx|�Z�ym��9'_��І���3I��cϤ���w?ܞ��]J����M�
���Qe���_Ld��
4���Ez���bc�rӓOW���q!�~?���+�;eL��o��!����a���-vӘU��]������Xt�1�Bn�Uy��hcsl���f��@�x?L�8�	6�|.~�O��O☑�oTN����4q��J��L)���ln�u����-��n>HFccO<��� }Cg,&\]���Q��:K3%��15��=e��o�
I�+�>kƐ9 7�P8����S%��F�hHd���rVX��~��>׶�2�_pH��e|�A^x��'�%�N��Pˍc�/ ��BF���2�O=k�㴖�هl���r�ʝK�(�Ө>����Ũ�$��Ů�Y�IH��H��;��lfT(�t�%�R!k_*}-�a~�U�Sv����3{�J	?�=6�%��e�U*c�oĞG�GR���T�v�=� 93�[_Y�jaL��VX(Ϲ���3^���=�����,_��h[�Ŵ�g`b�kE<1���m,�g|�vy�E�*0�;/8o���������=�n�!'*�<1����#w��vjӆ��ۗ6���p*� Ã�tQ�g��z�Ѓw���U�_�}�D�{~�c큶���8�piy��p����y�N���p�����4�F��f�\'�e�X��:�v�[E"�.A�\�O���D.�|f��yn��/Z���#B=W�A.X���q+d�?܅��G�4m�'���BIU/�? 
C��R4;��Ư��4F<)�cB����"�qD�' �{�y��K��Sj��J}1�]����v�҂��M�W�����������$�U�O!��8XcYU�
�M�|���R�+��i�8(Z8�%>�)t�rj kdZ:�k�j�85����F�+��
�؅n�`���+��U���hM=ź�g����Q=%�?/������0#G��O�;϶�v
<A.�gNJJz�i�S,q)y�d֜X5k�w�����m<4j+�B�.  jZ�iLF+RuU��qa6�)�%�����ۓ���_��5h�J��c�dA��X1D.Ν4�S6C���w��%���G�	i��c�"wvw��ގ=�ʝ�Z�"�͚`�	NPd�`4�>�����=SЍMT+�[ЍpY���E�˂���:�t?x?*��->��%��6ÌY_m52�i(��	l�x~��NT1M�k�J��	��W��$�G����ShP^�/e�_�~�#��J��c�g�?h��`3���Xa�'/+���e6��z1b�$��xf��g��,��~TX�'Ϧ�_^����Pʫ�ڌ)bcvr1���c �1�>���M��؛��	[��6�z!ĭO�N�v����Ԁ�=�##	��s\��Tܵ���$Ƒm&9:.�a�#B������l��L��t+��ϑC'X;r��s��S�m��$w� ����~���m�r6���������E��$�őb
Ǽ �$�`5�z���ׁO�� �������Mf���ĳw�
�1w��]e�j֌�
�@w�O�)�����:
��.}
���9��/�1}(]��|��
���z=��`Hf��<��%
Q5#]�������Y�G����S�t���:��%2V��y f����h@�ݫ���/�sGp��r޳��m�g��#C���n�|λWN���4d!euќ�9]םd��Fû�Q���{~~���t���q�gަ��(c'�R�4_��9���L�:Z2�ּk���lI����ug`��b�S�YJ�1 �