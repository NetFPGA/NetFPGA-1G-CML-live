XlxV64EB    2d4b     a80Qmcz.��5ΑW�T6�ā�)��ԐZ�E8�չ�g'π���z�^k1Z��3���}˧�@Q�4+���|4����>�!c[=�Z����h6N-S�1���H�m4xq��W��Ӊ���5����d�[X0d[Ε����x
� �B��b�qp����<�Abػ�p�[�����T�pd�㣻I9O&��`��kj/^���{j�>W}�.�=�N�{�Q�
���x�����ϐ�e�/��p�^��ⓢ/e�D^D�����=Cr�^��!UҼ��^K�E����b?v����׹_����kY-�L�o��;���#�)w�.G��,���C6��Tp�V����)�Ym�P�œ\��t�"��a�b�e oo���q��
�Q��_'��i레m2����� B+;��
w-�4J������1a���7C�#��f"���EI��,>q��� �m��ک�/���h���A:;��01#�S�3}���r�#�P�tWQ��|��Ey�D(�aQ��Jf��T��0ݾ8�{Zm6Sߪ�Yp=���L]�"��5˜t]j��f���& VвPu�:63���gL��
�l>�paڳ�rw�;0eG0��N2�?��l*�%�����u���@W+�t$���Q^D�or�GF�9xs�֖J[T��J&���Hз�|κ��E��8C�/U(T;��$(X�|N����125s	�|3�7�,� ��&��Lg�|����V<�4U@�W�w���,Ķ
�[�?�X��+� �d���_Z���6�`�"A�[ŀ��s��w<AP����6ua�L�!%[��Q�c������6��<Б�Hg
� V������V���u�>
k*�=|��t�xfM�k�Xـ
5��AdLqGԗ X��o��pP9j�i|���m�$DB�[�M�*���B�5N�³GoI3 ,㔸�π���+�[B�Է��$��R�o�:K���rw��ma�5��zk9Y-4�-D�g�-� ��6r�s�>E+��q���5�ڭG>��f�`?ӍX�UNg��DD��V_\�s�� &T�:�I�X�k��3?gaD߼)�_�2js>: �]u��� j4)�.���hĢd�Ů���@�@BT �Ei��񳍕H'�:�`
2�LQ��&n�������Uk� G%�A� ��{Dg��53��-�:G0�S��|�2YK�܎�1]p�m��}>9�t���q��3�ݽ�QOKc�o��]����J>,Pc���q)w,J%��P�5S�:ӒP=g�.��Ha0��A�a*�K��E��`�!�ޓ�%[���5_A��j��FS٭�-�4'F�C#�����&|�N���T0� �s�V�$3$B�ñ>��Ⱥ֤��*ɞR�O{i����/�%#��8*a��2��L�R�9�!MBe��^%/悎�8��*1MP�N��)j,���IK^;B�2��>D])�G��n�4xaU&�㒭xŜ�thY��zY�5�Ͱ�Z����&�+�~��V�J���%#��u�LgZ�3����i��K n}c��I$�l��:T�2M>��<aΣQ��:�FtNc��w�F�a^�]���qg��m��J����e$��ۃE��ǧշ��$T��Y� Ɔ��}qg޷gR'@�9��ۭ���>v�����w�̥"(�-?Vӷ�&�9���ʃ䥡��;�zn�K� ��(؁90Ё��6��)�e��K"QS_iij�)J�bЧ)�`�Ja
	�"4��l>cւ���^t�U8�+�_M��^0��
t�+b|O����J�Ǉ���}0�X�ˡ�J
��r����w[�߾�#s&Tc�[�3;����}[�AF-=,p��}�G/;o p����X�v����U�F�z�&MF'a>.GU,q�: YI�6J�0ķ�)&����:<U%��T�q s���ȦJ��,�YZ[�Jv"M�c�w��x��W��`B	�4^×��pʥ�]j�߅�(����!_��0ܝ>զ�K�nۖ��M���R�h
�4�lg6lZ�V�F��l;��_��ȼ�����L�� ���s�3\�`�P_T�rQˣXb�?��A�C�3�`n.�&<U��c2�ob@�\�?l�sBs�#^�_P}bd�̈�bM3�N�7"���-?�t:�Z��񮫴�Fr�rꆏz`ϳM�u��%>4E*�d-��O�'I��]�3���V�v��,3��˔�9�|F3�l}���beR|����<1|�XlP��nb�TĔ��ә_��e���[��8]�WZ�,f�&=
���Έ�P^�QN�v#�_4�)�^�Z1�8�q�7�IM���������n����YK<т*)E�ͧ���g�!�;{�NN�"��J���z��uR�2���}�a"�@!"�Ҳӑo��{tZ�QTZ����<��^D�a&��q���{Ak�EB�~�ɧ"i��;��M�����N'W��`��'Sv�C���}O���韫�	�� �.~R��,9ӷp��Iۙ;�p�Ǐ,]�z{�/��Zs�k	{x7��������5<�Q+���gf�G��(*��8o��s�r�mw@����;�o1�銛F ��6ڵh`�["S��}��ֶZ�����.8=�p��z��-%#���