XlxV64EB    39d7     f10H�Z�jg�iܞ���X�2�UJ�)Jp��$zx�K_~)K\~�{���`�+M{�:�&������ �y�q`=���;$HI��������?එ�/�N��>�B�}�/n�N�sd�м�j�/zhbw�8�P.�A3��^Wz�&�F!��o mY�-A
�+�S��cu�S�bZ�ё�?���������{��+c`[6�JD:���uU�Cr��3|0J
��{c+�A�NV������Bk��/�!����GA|3�]�G���"�� ����YR�y��|�#�o(id�>K*� ]��Oa�| ���i�A�������<��b/,V_m}���-�uUĘ��kF�i3��܋�^.�ӣ��L���83I(,Ŕ�/ox]JD�B�v�hT��H��M�ԢVΔ/|�� �X?r����DN��G�+�a�v0MB¦���\]1��V�C���u�Q̡,�_���'ð�P��֊S�s���?!۬�6�|�����o��uP�Ӭ����6	��U��N�Ëg��v k�@v>�]���w�����g�"8*B��C"Y���@-xi��r�6Gpj8�#ʠ�w��	:�a��,V����9������(���e��@��'�Փ�n���˩I��#Vz��K�h��&iDM=�)�I?���}Kݼ�ʺ�0wQ��,��eeAoaIe��3��u�I�+���%K��\jv��絻H0hDo��&T�و���} ��;+c+�8w����9%��������?${t�A>G�V�osw���͵�h/T¬W2Um�؜T��=��p�)��y�JY��dh&��9���Fy���P���	x������'_o2*�*=;�ǥ�?l_[�s�d�Ob ��E0;Zl+��7Ml�Q�k;�Q�)ΪR7���WQ�������s��a����"tL@�N:Ǻ_�_�usӸ<ź6;uY՝U���Xµwaų� } � <��ʹ$�����1^~�Je=���6꒬v�w�$�8��$��(*v8�x���j��!pp�nA�,�;3a�Hu��������ĸ_6�*D�������|��YC�'��k[�FD�`Q���i?=�x��f�GL�i!qr���e�}���u��ټaat�L
~�jr��#�d^�?[+.��PZU/�pr{=�Y�֕�!ڤz蒐n�r�X����)QQf ����EP&��.���ߍ$�;��n¾��rY)����DI���^wu2)~��G	ht;S�5����Pà�i�)4�X]mr��;ܾy�m�	��'�1��e�wY6���	�T]����9�̆�қL��X8 �G��`�褤k�6��V	W��$���\�W���i���A�F��~�܃�"�]���_|�!\����=^@��7��*Z���g
�n
hEQ�w�r��;gͱ꛷��:�t�Ѿs;(�(7�(���&XT�X�Y�/�֠P�!$sU��8���;�g�������[hU颵 ���k�΋$��҆娾%����NY򭯺�ZVp�2����N�mso(�I�l�8�ѧ���Ⱦܒg�{�O4��� _#�@NX�KJ��Q�2����'���/���EMg�ev��� vm�I���xsN�JP��������芏1����~N�mGV�~����D�䐨\��E��Ӭ��Ӈ>E���s{�Ug�`���Y�M�pv���@�8�}뾧L�A l�+k�t j4�
���p;��6��e��5(/��� ��"4���uE�bp��l5Ђ{��+
����|�Z��Q����e�n���m�ʓ5ek�L�I�¿����#�g���� ��*{�B.D�[|���>�=7əv�`��AC�������ǹStZ8*#>;q��a�hJg��-��j�T|.��U]1?m�C�LU�.N��d��˅z;�6͹o�6$&��N�K��f)�o��Q�h!�D���82��Td�0Ut�4؂.��i;�!����<?��pֹh�>��;	�
6�Ph������XU��54~r>�/�J!~q���g���T��"���g�ҔhM7 ��L���
��
�M�T6�����ZD4ܒ{��~������U��
�f���y(-��G�b:�WӃ�7�H��*|��>X���"��)/e�9����$�ãVo���6`<����Χ|����aߪ�[2�&wb�f���C��L�����l��L~�d%���Qx��zS1`��9>P;
L��#�%k��hXz$��ZV�����~�@��.�=�|E(4W�6+ԛ�:�G��� $VB9u�Ģ��o���Sj��H�ٿ�H�Gdn@r�f�o�~�����	C"%k��Ac'�^�O�H�	@��_]8��)؄+N��*3�"k�6>���8�� %�������j�{�<�-����W���h�N��`�۷ݪ��#���h1��鸔q_����m����PHiN����Ji�z�4Y����j��e����U�|�^P�#BH���ɱ۝��zx Tw�;��B!�%�d��v�CVK��~��@=�f�`�9�Śѵ�xI,��/<�EI�}�[��6}f{���]U)�~��J�A4bz� ���y�����f�?3�=��E�\ʥ+?�R��u��u���T�����R������$��~�1sa e*<<���ZVq����fC�V��r3�8z 6[z���?��g3� �*&�ՑUУG�$TQT��ڕ��"tԪ/������Y��tF��qS���{�n��,u���W�7��˳�H�g�3����a{�}� �N�>���ӌ�����!߮c}ν�1�o��A�QJ����bH�73J�-����ʰ?��%�LG�TI���rR4$ n��ՠ�/�N��{n��y��T=�R���`������Af�KQ��u]�:0gsC�"������4�Hek���(������y�hU/htc$SX.;������-Yy������b�/uЌ8�H���:TY.�˧�R�Ce��'�>�T�� ;����)�frf�Y(�)m;g#�����Dcs��kK�2��y4������z�Ǽ1��U7ŭC�te�h�#�YT�:~����m4�z)������p�:�'�ul���B�yY	gqI�*��(����`i	�X������������J~L�.c�æ����5b�^M����_@A�¢a�+{f_e�����&�5ֹ��΄��M�y��Q�l'&���r��N�$�2�?3�]��?�R��iC� e�ԿD��| ��N��3�ڷ|žؓ�q������]�1.��6�	Bʡos��nI>RGx:�n�kg�\WN�b���]��r�j��'�I1���!rT�c�\�tj�ydP���J��<oq@��D9�O�3]~�p�M�6U�)~FJ�<ٗR�һiY?���%n��P�H������&4�2���L}�\�*�O��:�X����{���)���r	�K}��w�:?־N�� 
�;�Rü >stNp���� ��t�=M��x$:H�y��ME:�T!�����k�E���W��vgĳ��q�=��J(��}PZ~gؕrQ�����+��ʧnc��_��q�Cމ��ls[�������[�>Zݟ,T5�2$\گ��QW]T���k*��Rf�L����Zo��٧[/��	ZހL��+@��؂�C�iq��U������#Cw�6�a��s�u(	Z4�� ��p��K�x����@��:��Ѩ��n���?�fa�� S�4&^