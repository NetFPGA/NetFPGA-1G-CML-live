XlxV64EB    f830    2c90aΎG���������&�N͑�ۻ'R����W�	�	5�.l'��\5�=���W��Kj`µh�I��eB�����՘�� 2>��e "�~5����yiD�L��cE�S�+N�-#�j�УT���l�s~�m�\�0]D�+;z�?\�;F"���$�%��?sL�n���.�Ù��ƱJW�*S�W�>��B���wa-٨]_e1�9!��g����� G*S_@e���[�5>���'D�K
6QE����_m�%4���-<��ԍ&�G3%�\�*��\��i����"_m]�ot�h�{�G+T�!z�[�����0�f&�X.y�k��\����i�w/���
�hs�`x*�3�\���!R���A��Ǽ�$0<�Ҝ�n
�'4y���-�;��W
d�j9��e�7�*�sgQ��H�E������ <�B�R&��З�\�|�ᜫ�J[������Q)��w�4-�-E���?��&�� �~ɈB"�]��L�K���]vˁ��&��l�	g��A�	ƌ�!��⃁�
��"�+P�l|Q�'7Mc�<wK��9���o�� ͢H��:�8n�G&b{���aT��������s	�2�?���uZ�3Q d�����\�씵��Y��n^7$xDX�"���e��Af]���n��0��F/���H�A�Ӌ�`���5E<\��Id���D�yʌu���s��ˢ �@?��=g0���>�����-_�����p@a��f($ҷ'������_�C���5�5+�d�9<��'&��?��r]�{\�{O�DA��8����_`3	&MA�}�Vc.4���.H�+Ab�~e��aC�;l5h�����*��]�����ե�/[�hYbD$ZY�a4@v+�$�K�k��ZS��6hpy4;����YV�4�Y�,�)}�]���]�d�W���t���X���ŅD���~��/I���\[�5��2Di�n4SPrejK�-Ȁ��_ɝe�$��Pc���C����AU�2�W���-�eƈ���`v�}�G'�3ĔD�t�*���
��S�`y�y�vIH�]F*�0k�]�lq\22�&&ؾ��8,�<}5&��}ɠ���*���>�
7B�Ŭ��3fJ\@��&d�=�N�+"Pr�{w¤�������H�IYq��@�TtJ�
Z��@�'A��Pխ����t��*'4U�ugM�鵌�xi�2�qa�$o�;��AO�sq���L}Cf�6�aC�0�j>E�Z�g�A�������0�<�UXم�7�����7�v��L���(+e����"��1QɅ&��W��<CM���
�]��x����׷�FN�Y�s��a�b!��(�;���	�M�*;��	��濆Lɏ�!��c�R���0P1��"��6w�z(�t�xu0���}Yn�#n
fsN��u�{?���/S���s\Ӿ\ ����=����2�� &����,�y̅ZK��$W�u�C[޷�̗�e?,>����H1�,�1&��g�W'��Yp�8h�6���'g>��%@4�{��wF�Fe�OѲ�)����3Q��2k:���!��r�aP���-m���>�9jk�\���v�X�@dCE�sOpK����B�Ό���C�b��ޟӼ�c:0v����g_A�i�)H,י�bST!�ĸQ`�7�i^NF6P�[�b_��);����
sja�{ ����H��	��_��0*��	�b� ,�m�*w�u�/��k�p�CD�PW�.�J&�x%��MI��A(ԂZ� �P�Nԯ����]`c���Ų����vH�V�^q[ds��H+7�.9� ΡT&�@{�X��H�F[�c�d���5�93���^��lO���( ~U�q���,젶�PF�w��m���H=OjL�[Un��s\ !�:d���'U K�fw=��h���u_Fo(I����3�Fm��yY78�t��1�J��	o�ŀ���-a{��a_�2����u��	 +4��z���a� �;��DV}d&�r��mM����,��A#;.qM�0�R�&	��eF�O�yG�aWMEӓ�Ťg��̅���06	N��h����Ow� � �Y�d���Kٖ9��ێ* a�I�A�����CɥOGd�@ /�V
��#���"����>�I��'�T��m^�m��ɖ���e:`n�R�t��X~�J���bZV_q�H����4�m@p��%�`FZ �ђuS���VN�hDsw���_�k%)�r�H��7���!)P�F���륛T�h@��3���hx7�}��@0��0��R��`��?@�c*��uq;�@����SNݎ������SO
��#�r� �j}�ЎD���d)M IT�㶷�Y6k��ԣ���H��3xz��פ "M[pT�<=���>az���q�)N�#&=���|���gӝ��zfu��q����7�!�*���Ͷ�1��	�/��X=M��p�����bId��Vx�0}1�u����s��Qtp�b���u�g� 7�����/.�@p;C�O�YZ�K�|9M�z3���~w�Z��(L�hZ�Nb
S�r�C���e��d�#BS��$hyv�У.t[H��f͢�����7G+��x��D�=���C�+�cR7$�;�Օ��u�Sa�V�Y!%?fw�P�?�L~n�����i����O���H)���g,?�y�pȤ���Զ�?g��!����j����}|��������$YgqQ浰Qց-��%t��QC�7E]߅qk��ζį���m����z�9�⾠$,����p׻���Y�Bg�����􃞨���*h�@MBhz�h��{�w���%̃�8�[�<�Ir|\��Am1i��,�%3���c���B�8",��ޤ����KA�Cϸ�s�$����&��(��e9�ө��ʩU<�E�q#�
���$Hp�qco��Vn�<47�Ǭ��^����.aͩ�2��6Iþ�!�jGB%n|�<�d8�	��.^�O��O@�,��ϰ�n�\��}k�_n�H��x0�]����$�<���(. �@�G��ϭ�:���h��)�OeN��'��]Aи������	~�x���S����a���}g����y3|��_����u��w��	U �1xm���H8�QmUMv�<�����a�%����[��⦸/�= ;�-�r�kn��L���Fʚ���$I�;0�GU'JX��/(����$?׍aIO�C�K�j�ED>L�����DW�����'����ݺ_Ș� �{�]qQ��
����2N����:��H]�E������������<�H��I��H�jI(^\29$v����A�d!�?%�螺F��`6\���j�C%��)i�����׃�z]s\��;�?�N���n�7�T�^),ѸeBnA���$R-�ᡌ#=:y���O��n�^ t��u�% V���9|8-Q�*�/�o�u�iT�����7[����W,eQ=�: �U2C9O��<����^$���e�w���sf�m�g��%���9����W�7Å��^��I���e���]�{gP����F_�����KX5�j���E�P�>l�KD�ܛ�B�d_���?3z�׶G�Ħ?0[�����b� V�J�_NTUcs�?�s�6f�g��>���d=5x{$��97m��)�6ޕ$���WD+l��ɮ���Jd�u�������B����;�)σ�*�1rFe��"H@��4 ��m��&U.s��kT���"6o�4��i��]��B�r ��^AP�����JJ�x<C+@��x�^��w�T1��� 4��|��{����J\���ja��+��O�O߄B�S���T��1�g�b���??5n&�peU0&Z=kܑ�sm-J�0)p�%�m�����y�-D��`�@�[� �Ӵ}��4��N6�|�4W}�0��h�D�v��S�A���|��~Тe��zl*� s�f3K��GQQN�h�^�:��Y>��54��~�������C��+��h�L1�X�i�$���/�n{���D����a�3o���D�*�-}c�x��_�l��!��^��� 6�	8��C����;=`�)�`����ĞNE��o��?t<�F��^��� D���bi�5�;�e�Gݥ)Y1��M�ֶ���-ķv�B�r{�aH�ֆzf߭D�*_����\�M��VLoVV��$nKw3w�q��N*l��5�9�����윗��08�[+ŨCY4F���[+7_���/��/�E�#��c0�P�eej���1�g����,cz�v8&~	�ֽ��'�f�[8��*^ԋ�g6�2��υ9��}�v�px���B"������F���B���/�c"��f�ҕcLS�c}��R�v�==�b��d
� ;�o����]Wul+kf�E?6�de �_��K*�m�Ŕ�{�|]��@zd2�πs��@sҎ�a��M�����nh4��F������s�LS�0/�gjy�� }Y���)�N魜�Ӹ���~�,� �v\��� �σ�����0�[z~~����Lu.F�%���!2��~ң㲚˴��:`{z�`�}[�Z��b�m��5���l���ĜjϦqLj�K~/�\�0�f��MABsD��
�����\( W"�#B��O��� ���Ѿ��W�*g�Rz m�tx�.���Ŀ���,�����'�P��	д*���7��7%w�}�S�3Z�x�T�82����5z�Mf�}��&��c�~ O�yLi<jf��~�x�&���84���F��*@��%����J��e/�<�XȀZ�)��nMU�`E5��&��@8�D��4��H��H��hԑk�|����ɦ�bHÑB��@���ײ>�am�!���X�t
hᜍ|1�2���؁%R.�Nx�����\���_v"���9&z��6�{�Z���.B��O�`�F"�\�@?h4�po��J�&K��Rf���rܩ#\��+E��pq�}b����$jmed������r6&�A�(D� L���ڛ�&�wԤn�'� ���B����^:�_b�F��,.Z/&L �z�*��t����S�,�����܃�H����h�NE��Ox�Nؽ�i%k7ϐ�cK��v܅�S ���{W(ފ��p4|[Qlj9��5w��1\ (#G�A��V�P�bp@ae�Ќw���D��]��2���.�"�UP�,Ű��]�WM)�>1+���Ch�I��_S���F=��  ���c�S��U2��$��9r��n��P�o�>����-U'y�>�=�q9��8�|��u�@Q�iB�Ȋ��B��H���Ń[�2�ޓW^�?VBl�Y��ie�tV�H�c�	�п�M��=��3��z�횩���ħf�x������`�)�h�ܥ�9�^qogF��>�,OX����IJr����)�U;��+���m�2!�ΐJ������puh����]�����l�t4���A�S�oQ2�������������[aR���k�;Ǟ#�M!B�ok��>^��8]�U�܆� 	k홟��f�i����M�zV�ou�n��W5���)t����j�׆Wu��h- Μ\J��\K��ǽ:��6z��
V;������8�@ZSa	Y![s��}q�b?��YB�CJ�6r)��.�س�/5�ĵ�y���p�}f]@�f�;�t3�92�M6M��� ��&s��%շ���r(l��4NM��d�%z(��I!�}2S���s�X�?�?bbj<����zo���u�0��P�A-Z��薣T-�?H^�4;��U:$G����W9|�H�ŷ�6�r��xXC�_;\H|��Q��1~�G�2��k���҈D��|d�D�\_m�6���v��duM2����}[?�|=�;i�����+����Ɇ��G�e|f^ۅ3�7���LptN��~�.��U�x'���-���C�R�f�!���^1V����N�)A�������� EH}i�,����*��S��Ϝ�ߐ��h�'�$��˼�-l��jZ��j�etr`)>b���+��M�P�Kc"�m��gJθ����,�H�;ɬnҸP9Q��,y�FAT�t�]�(T�;�3(����Oi~�+~&4S.�����Ad������ҟj��u
D�B���.�3�$�shY�S��q+� �p�	��#�R�3kx7��XS�\`�"-����gZΓ��EƉ�h`]_��sϭx7��C���?��:_��3o��e������g���y��yE�3v�������p��`K����=�,�*�f��vJ5J���%��_F�E=PZ���A7�wf@�
��Zr�v?ml�3����#��-�HE���͝�NS����_����gD��6�O�be.�7�L)"%�����|պ`�W��Н��J�͹�ě�+�ry��#׎�V媫�\n-FȂD��|�'PJ�0Jz��'�F��x�N\��3.��w�Y�����Fj��A^���^�UԷ31��eo=�f8�o�c�kn���`��<�;��ڦ�d�v �3��*Z��|L�K��x���_�q�t⚀��!|8l��HA�d�M���N�/�^M,��2�����$T�m�!�x&t�vۻ���X�x��|�o�]�M�߫/�G�/�w	��g���3a%��g�\P��cA(0׾|�
�l�w�����lC*@:��0�����]~t��~;�5��T����=�����]�)#�S5��8@ň&+']�YĚ���\P�E��9���j��P��e@'YH�l���p�XNo����Z�t_bԴҫnoƽ&��Eك�(c��w��#J���"A~���t?�3超m�ɦd���:+4\��+u��ӣ!�sH���AT|���P�f�Y?d�E)=�A��f�T��2V1�5��~u�8�8*���OQ��Br{�9�cv�f�X�i�;���XG��+�Q���b#^~�[�O
��U�.0D`i�_r�;e�36�Nn8<�ag��mm�e�]Vosp���rz��U P=~]ӆ�����Mq�C�O�i���G5*9{b�Y�=Z�5��on
�$�=���RW�wq��/��̋��v��j�E�J��x��r�;���+�̸w]r0�sG��>��lΩ����ThJ꾃��⋳�߀� _�D!����oC���� ��sSRڨ�i��i�=�3���!��.Y��T=���/�[^��SEDX�r}:!���ɖ�����1��2׏�A�8�2���:�p��rL�\^�o]p�$vT(�&";��m�Yi[%�����rGΰ6q�j ��Y��[C���W��i�F���h*`u��dE�>������-��O��!΍Ŵwt��!���v���)GԹ:ә��Y�!��MU��Pқ�N(�AH�i�^ͦ�����!z�鄭C�#}���u�I�v�չm�}-MB�14��]1te3r�|�͂4�B�.V��~�� �HQ�t|?��I�>~��3�'�>3��!��;�ڶ0^��mW,�Q�9ժ�9�N���-oecO�����Ǎ4m�-k����#*��?�h��pl��c��e���P��B[*��Z��S+�R�2J[��A�Y�ŊG���+
X�h�~(�gLd��kvRЛ���i�əQ��ä��sT�C0������y��u�<�)�{��+M�Hҕ4,�&�{����3�bSU'�و[��V/�^�>k�d�Wch���u����oE�3;q�<*�,��:G�R"�r�8���o���~M�*%+���C66�F!7=yy���O;�b���C��q]��J�ɚ�X%Wa<(���ϰ�n;��#��� ��v��4`2�SΈ��m������[~v2�Ů��V̚C2P˔�w}Tp�@��c�Y�m�$-��2��~�9d0KaUGC�I�e.��fªg�'��̈́�jp���ǁ��.�����KH��!
 k],�Ca���*�.]�ັ�8쒽��H���1]��$�e$Ԯ�j������_`x��tq���F��C|�6���k��n����y=�=�\O�
-!�eF�A:�2��?�0�u�P1_�+����	�IH�Xh
m:"�q`��h��e�-��:�Z@D.�#�#��,�2��uFy�"�����ůE�������T�?���K����&Y�y�}~����5���Υ{1i}��o�7�d)�_▫�X qs�M�4HTb��U9�@��X�!o�,�x��nFda�R������dr�	�����Ҏ9i���}�j�މ��jΛ�j�2涳��AYYE|�O�w�߄X_$��� ��"���W���}c���/h7ي�d)_�ElqE��޴4�G��V�&���=��K�qB��s�����
Gw�Ph'���~0�<'��w.Ƃ��蜊0�����4�s�ز.x��57�m��%�i�h�`�W}5ق�M��e�g�z�fm�xoa!�(;��/5;�&�����{�>��w\=�CA��t���wj�߶�������F���0�Rkǚ�C�+�T �j�1J�\�Է^��!ĝC��^�x�����A6��V�AWs�ϥ�w�.���Y�B�؏��!A��
_NN�ᄑ�<�EB��pT"�H�e���B`Am��22�v�h[�nP%�Y�!�b�>nT�V>S�6'�?ڀӈ��zjz��0��YS�/�<���dlW�i׬n���%��BR��0��%d��*=�g�тѲ'̉�;�����������\.?1-�l�����Uu(�8A�Ǣ���5��d��r H�6��G9�a���Ii}�z
�n��V��d�Ϫz�*!aG[#�*�;�����)L( �ٰø��H!��J�1<�%Ξ{nϼ �j�
����I1��cцqdH��f����A�LZ�W� ���aG�Oxl�Q��J���QU�!�Yr ��Lg�|�gr��<$���b"������������J I�t+�7S�ɓB�~����-Ԋ����4�~ i�^�)��Vn�tOv����T�{K#���}D5�IA�p4]��g��v�U���R9�~J��6Q�eX7������@���V������ZS�$�xz�z��7q�5=��U�ctb>��L+�ee��/� _Z���J0�ecoU�58�3�_��p�Y��v|�?�>ڗ.x{���T�a^F�v�E����Zd���v6��v~pa��JD��><�?ͭ&���s���\�f���цQ��奢�o��i�݌����":KU��T�������ywF)?��ϧ}�ɒ�_�Ljد�1�v���Z�,'�x;��O"�����L5Uy�4����N��sqtx���&-M$n:X���r���vs�������G�[��/osF���f���$���:�I��%��VhT�3��� :FiSI�3dc�/֖m�~B�>��G���P��.���il�(�[q�M�.B�ׁy�%n�K�bD�>56j�<geL#��ߖ�}�E�P���d�m&������D�5|C��z[�ṇ�37�:}o�  	��3�o�dc0�F��݅2��y沗	G`+�/����7\��n�
;
�`'��+�� �u�7�:~�oU��Tr�E-����ބ6!h{�*���g	�Y*]�u}���$e}99�' m6�!�q߈�P��p!t�g�?��*c�aV�{����=�&d|�̤pQ�}�9/�M��� Ĺ�����џ�68���B<	ۈ!(�Z��6��d.]�W����޴t��a���� �
�O�	}��矹�Zc��B_��6�����F~(��2-�9h��G�~/M��*�[�6��>�������.X	�m0N�C�DB'*���	N��Tv���|_3͇me�n���EP�GmA�u��X�;��f2��av��TA��8���
�>���i��/����[���͏:=��p�ߐR������<��峋]H.���w�Bf���Qh{L�*o[8���ޞ�XG�?�j�|WO.��$o����K���;H���dc�����'�_B���Kb�j;�ձ��	J	�����]�`�e�*�3�;v�v�clʡ?���{�Hޭ��]z��7/ӌ��847 �Ov{�l���Ny+1��G�[�.�����kU8P��%; �=<Z�*y�h%���\��|ueQ��e\nZAOx�eW���D�9d�%|����)$�KW<'w7|��'��|c������7�9�|:K�za�k�����.�P����4K-}�qǨ�l��viƴk��Iٙ�ߺ�XdR�՗m�M������e�7�O��q��0:k��_7��zc�P�Z<����<���8J5���t�j��D���H�K�_��	5ȳ\�w����y9\5%d�W@l�1�p8��i&�ݝ���I-�Zhy[��'u3��;�Ķ�!��|eŁ���=UW��3g�p��h0wP����r<t�`�k�am@��3XZN��/�6�nyz�������k�Et?-Eq~AެD�qc�ʗ���v���$^)x��0���s�����5��U#����i;�����=��������z쟞?�T��PҤ�.�������)G�#��#��I��1�!��X4�w�J{�R�K�������i��-���\�-h*H�NS��� i`�3}Td����Aԇ:�ѧI����K�BC\������Et�5��{�����uL�������\#o-Mb@�4u�E�}�$-TP��=��q��R�o�x��k��4,����t���k{���|q������c�Sujv��n.^�nAo�6�����h���ϳ�B�uYNӕ^8i�3��0�!Q׫��+�(��Qԓb"�:��BW��L�f�>?ń��U�I� ��Bs�nZjHװ�H�xY�.����c�=;�q���	��l�jЖӋ�{3�,����Q��ip��}���ǳ��@�4PcٔX�w>;�G1��so��0tKc߱�����Td��kKR�OpE{���\�`�g�Z&�肐K�F��Ϥ���T9�"3
�1z�	���*���"5��O׫�z��4��*�� r2���ڊ��