XlxV64EB    2283     b10HcxF �]\5Bm)��(^]\?� (���RL[ ���(�>6_)SS$��J��Q	���*��!|���e۾�F�!���aM:.g�:}T�����$���Ɋ|�)��j9�r�e��<s�Y��;Z�VLK�8�����Pa�Hy��*�TfY
�~+�/`H�J���N��׸��Q�L��~E@�ɴ��҈��F�h��l�C�E�d����Hg0�K�� �IŵP�b2p�uqA�a0��.�a%c��(�ܪ&�y0�kG�f5)��|���T��11E5�($��nS�S��e�ޓ�h�֑-������a]�{}Ҙ{��t�����=��m�2��O����+kM#u}���U���}��?��I:U~�f�M����M�Z�c���D�[H:���3��-�x�X��G��h
27��G���̠f~2�O�K_m1`��{���=i�����1��V^����-nV��S�}�)�8�.qGT��.6�OLu��_wg�ġ)b��w��~bA�;u�,�x�8#A~�~ґ��W���{�;���Z)����=�� �܉�l\=i߮7�W>�Ձ���%�E�4��%��SC�?^��� ���]�bZXI � 7�� 7'�{�i��o/u�<�w��r�e�f�gỹZy�j�OR>�bm{yF�{��4�|ı�0&m���X֨�9@I������qu$ ��V���{�4W�[*�`�s�Kf����-�j	�U_��\`Iym6Pq��Y�d{���Z�Ӝ;���oV�d��������&/[�V���4ܓ�b�Z��������?W��_"^2�����庹^�3,q��*�HJ\
`2�_G�.�Z)��g\�tJ�B���	�ڴc(�ȱ|r�4�D�~�d�`tQH��5�s�|9�#8�X�����U�ԓk���:&3˻:�QUV3+3��ų�i
� �MVY�b/!�DЦ.�#JEsi��;�5��"�y0�����l�����m���wL�pF�-�	^��M�U�L�
��3 ͵m)3
d
�09�=��:W-3X���!A�n2?
q�Ƴ�@�����t�S�be� y�#��0q��\�l���o��� B�y.4q�=�_g���}-Tkø4n`^�R��UzWdeL�w��桇"�{���|��p��H|@a��Sȋ��q����$��[SbJi��ݢ���V��������s��kRX9��of��z�J�ͱ�+�|�JDՠ��<A���A�oIۯ)��s~��S����iP��!]���T�����h�8��V�	,��C2�UT~�����D�EA�n�S}.dG�w��A�XI�ҷ�H�՘� ��~$$ ̌��7صHu)��!�f2�lXO8���ˢ�I�ݸ��1"��pǥ�8
l����[m���f'��V������~X�v��o0�[��ǰ뒬�k����5�}SJ=��k�+���`"����m�e}�|��e,G$��׋L"�㖠�
��O���L���Ih\
H�J3��E#%����fdC׏�܇.�#�R�}g�gՁ�d�|?�s�RB�����P�l�IP�mT�5J8��ס��x��״W��3N?��aA��9����՝���mˌ@�H
lwy�oi�8i�v��G��@9)�N��6�SD�H @G$��6��ԆK�=����E��a>)�>w�̫�gID�,�rU>����G�4�UA;O�|X�F�SH�s��1=!������5�(�5������yx�����z�3Rh��gk��h@e�H�z��I	jx�TQ⚃q�>����h�Q��VfL�,�B���ܘ
A�:oٕ	�ڪl	c;q.�cb.O��� ���U���t{��7� �]������U<q���j�)�`9w��̟���68@׃ �l�Y�b�$�\��ҴT�Q���7�̊b�2n�SI+ȟ�6fs���C�(�
Y��#�]w�es�W�7*�^B����>=�̆�;�������_�z������nH?�X�Sn��2q8`6n��"�鯅�h�]����nq�Ę$j}�f�,���x(T���ƴ�=�PC[����j�V�z���֫O��`/��@g�h^�>I���Ѝ�+t�������$,�f�J7�W�Op��i�v��@:���j�^�3��1�*b�9J*�g�3��q��HU��Tr�~���B/m��I֛v��r>l�E]S���}Q;H60�3�Q��=��[Ps�䰉�b�R�	��d���-����fJ��S����"L�|w6xg�Aq�ݗΰD2��ȶ���{E��2e�=�״�q����D��ϻ}�B��r��p�Jz������J���� �u���s~�4h`�yEWQ��� U�.�HS�
�`�o�V�f~/SW����+�����imq[G�i�������|?	�VX��?#�r�W���htβ���Jg������,��qRt%����4�qH�V�������*EYQ܍v�ɛ��u
Uɋ�C��zR���P�rF�3q��V�N���s�K��ܪ���J-�?TX�=Et7:W2����>z�<m��{q#���z2g$E�m�@�I5���a�q{=�V!����/��.�Ciu�X�]l��&������]�!3}=�x�k�Pm��d��ܗ�!x'��/��9�7�bpr�̡��F
F�Ncr�����p#���䗈ۦo���!��:n&\��� �c;��Q"�;��!6����7ǂ,�se]6�h���$3^���&��wi�3