XlxV64EB    1727     870�̞g�Q�MlP�w!o���0u���4���=���جh���!����[�,`�p9������=H4�5{�M�
�,�<N g%��� �7/�B�}8��(#��J�<yU����g���M��UN�{w��j_m>|�D��zt�y� i`��K	�R�����c����O&C������ժ:����TQˣ>��j�A�����*O����٨�ڡ���'��0��*p;Avi�8_l�Ю(�n֤@bc�\�����ղ~�F�@�����*�nk#���SmJ>L~��h�
n�!���lh@m���3������݂��qTL�����s|��(Uq�zgG�d��p^�U|����lt]�M<���咜�ud�V��Qw��1�+&�NɈ�A~��^'��Q�wXXv�.�����'W(��@1,�|��)ʗ��S�xP�$����z<^݂�e�拨΋�;�հTY2Ӂŧ�Q�yD��m�C��E�*{���$>\t�S�5����>�9��g���$*_C��p���V�� ��Rk$��}���u�'a�ۈ����(�Iw`�1�%˛t�\�Q��_��L�ڥ2V	�w��dJ5+���FC��1|t K}�����4ZWs�	O��Ww��3^��åX���� x}R��Z��P?�:�eL�I
��$N��BP�Ȉ=,����p��m.D�;Q}�Bɔ-���a��b����t$�v)��CY6؛:z&����k�ٻ���y����pr��gf��)i�cl��@T�8��������).V�e�tŷnQ�� �+Le7�g1��Dg��s�� Vݎ䄩�cV(�W���8��%B0V��cۯt�J<�o���V�hf�٥�3ډ�x�c�/y�\�aLj�y��妚I�ݳ�k'�ښ�A,��rWˎm;��.�60����M��k�_H�:cq���sF���,�E�6�V6	�T~=��%�x��t����.8K� ��2b5LY	����-��3��i��oN���4s�Ġ.ez,r �94������-�������ѣ��Ώ�0�� 1�;U�[�p逘�2F�X�7�8�8���0	ܿ�*˔Ӑ�vv� f?����I��2=A��K�M� '6:�vd� 0A����Q����5�Pj]�#]��)[�m���������͹���7lz�0�MF������J�Ӡ�-��X6����������l@�����gfw�'��G0���2��K<*�BmJ��#�%#�<�/�E�;E�g�Fg��	�L	�����knq�[�ǳ]��A(�hU������luu����Z[�I<���"/'����;�
��b,|�|��������d�~������
ܛ��YA�I�Ժ�����n����f��V�"H�Z��dq�wH�M���}G�"ە�`�O�k
�%]�<�:��^�7Q�K�A˼���P��i�㢴|pѝJ���v��sm��b�g��=��S"4��(~�{G�?I�4�VFŸww����;~D���"��b�7���g kͯ�>��u���ڑ'�����<s�0}�6&�f���ZccS��ګ#�D�9 ��$Ԭ)K|(1�;Hj�a��!B%$���
86�N��W����^ꖳ�h`q-�8Z��*��j��:����OS���=u����c�� �RF+DX��R�R8�לs��)Aӫ����Jg�:����#{�9��niПmO�o��#_�T�-�
�De��&ȅ�3�`���/�X&��q�b�F"0�	�����i�ٟ0
��K���H��Ud��:��#�����#�"�*��	K�AV4�!��"<Ź̻��-��<�:�Y�(�ﰫI��J���=���U�K�ن7����>�~S�qWS�6�_���l�t:�{�" �=����E�{aw��X��5!)��5(����4|0:$9Y�:�j=r���40�k��N
���JiJ��mc�7��Bֿ��2.QK�S�x1�^v<}č��J�a��g����M�D�!�"��|�+��`�:��'C�����p�#> w���9Y���
˸�����)�8�ծG�{���5�ý��