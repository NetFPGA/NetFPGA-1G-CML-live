XlxV64EB    5774    1440�˘�G�5?�E7��qј�
�D���i�Y��Ǣ3!��8|㠏�bJ|�uZ	ר�*��ŧuq�Ћ��h��;)��?D�xK�[���3=�"��M�.A�P޶��'��0˻K��.�������F��W�� 냄�2���ּ��K6/��%xj�Y/K�i����J�p�(���DJ���!%�	;�2���?G�Le��[\�� ��3���-��@�c��!o��M%-�K���R#4�]R�@t@�׳��RM�<g�$Me-�:*��)-4��毬�eμ�#\��3�"^m�����ऍ���̤�</��W1�勜tS���Y&GI�b�y
�և�@��F���!�D;]�G ���91�DK��<���S�J7GV)o����+2���\�Z�g�]�D��B�8���=4��	9^�q�W��H�4� �K��ЍЉ�'2�"q��`�$���L���������W�y� +H��g�}��0��꣛��^�5P:� i��7�|��cC|�Tӑe��I2)���~��+�'���qX�hMe��w�)���+���h�G��Q��&i���
E�ȣ7<�vA�$�Ji��|��Շw�s�3�Ug�,J�g+�hwU-(��J�!\,XS�|���F)}oM22Ç���8h���2��c�� ǌ�X�'=�o�0.�� H�O;8"�������I�?��4 �*���� t^P�ޙ.k �~0ax*���}�o���(��$����)����7~�#�U�J�/�7)�������0[�P1��o�:҆�K��;��R�w����ڣ#�	O�Ȕg���ÙU�����|#��;��R�5�<���0�Tp����G~�]�%$ȇQ��N��p��;������Y>��4�`��>ڗ�orphR����U��q��n�Md��]����8tP��4@4��w�QHg�&u���2.��G�@\w|�$�C�?~��;��m&6�f�&G���x�9�9�ֵ\��Nז�I��P�#z'�����?82ݗz+�G9�\6=TQ�ـ3؅a�6:��"%����G�����鼿Ar�>ҭلj�����ɛd�����OǤi��O�<e3!��%g1�� /ڶ[t��.i��_�?��Ə��ҩ���UJ���"
�q��g\۪ �S8�B��	�_b<�pl�����K�0|>4g���/y��cތ&���G$�S�L����h��_a�,��[2���oC��a��*�Vx�~�!`Iw�X��Zcg�s+�e�)�H�к;5���&�(�sM6�p&ּ��@�G:��G�ݳ�\��(�eN��}�Fy��>��Fu��*�N��p4 �6�n(6]�~x(1�*]X�Cs�IN�ď]h��5�=�u��fU�|?��]�Ϸ	�SZ�f%� ��)�(���S��m�·!B��A(��9B9����;���d�N	Ne,M+�'i�E9z�?	X�೭��
�Q������Y��Q�S�?ϧ�Guc�>�NO�k���N��B\*���U�d�M ��i��uA7礄�R�l�c{y}��A�:|Q
�h��/�61����� ]v3���n{2`I��6h�a��lA/�H�A���@�\��?�e���̸K#K�����\u��<��t�ř��Lq�'��B��p7�MQ0ۓ>ιȡvW�G##�8��M��Q*D�en<�ju��ցt���9B�:M� �=i���k�3����?�2�������]�&����n������t��m �߹jt3�`�<�ꏄQ֕��
�>�(�6�k ��g2��P'F��x���x�N.~�1���s䨪W�e.���\\|�s�5�]�e�����Yt���Z���3�D��RV�D=6�:�W�2��$��nS@������ω���+��8�L,��'��˲G�j4�en�I	�g�`�.�pkѠ�GRr�D#�@��y
� xOM, �?��o$F�!�M:}W;�: OR��K�����K3!(x{I'"���:�P�!��A�ϐ�����}�=��$ɒ�T�#
���huhЀ��SbG�����Y-��w���[�X���N�Kx�y3:�1��4˨��@����$�%cgKAVZ����nN�Q�=�Օ���V�3L׆/!�(a�p���T�g$���o���'Պ��G<Qi!8��{Q�2/�J�@�����}?{�}����bC]XО��&t����S�	��l��"c��u<��� 
d��
����&�bn9��y���^P,>ԡQs:��ٹk�w~-ك����܈�Q��EC��P�(��N��,,q+�r��k�Ϗ� @�(��i_���7F���l�+��1;l,>��Y2�f4��1s���N������G�Q�Q��L@�w�����@�s�������01�;k'�-@A:S�I�b}PVs1:GC���D��22;���+�JѢ�ƨ��z�H�����k�[uk�1���9˾�q^���R����N,�:�U"h��|k����nF�Á�S3;�9ɴ�cl�P:~��8vb��Ö��إԶ9�~����Y�>S���g��ܧHi���:�4h|uD?|�k9�#���{��х��-�����o��vG��}�I:����,�|��V���l/���&�5�N,w��e�P�s����<e��ӻÝ����A�,۷kݖ[�}�]H���^��?ۤ��'(+��T�~���X��a^a���}�e
�;=��W�L_�+�}ד>gL�1�^���A���@�}Xܧ~(6��`������Z�Ft�d+i�����4���n�T�$D�*>����($��f�0�r��8��d��mt{�Jq���34���em���Pfc3���{�ŹO0>	�N�	��|�8d)\����.L�?H@�s^9Dj���=��l�y13�neg+"����m��� q�O+�f�M��KvG]�2��UaQ���{�u��م~�lM�^�د[��6p>dPu+`-���y��3�^����|f{��Ƶ�_[��-��G�sJ�"}���⺷=>�� ��S#���p�+a�ۄ2��c�2�s��u�>��G3�B��FVc@Ж$ԩ��=��;l\�ٺ���X3D���V��]�t?.���/$�O�H�����C�-gL�M_�1�aL�Gv��c �:�.S���_��ك��T�gn�qo�g�B�!��D	Y��t#����_U��h;f�������hs�y�GO{J�T�����%��n�����o�u@�	�����
N���`L�/��^RI��
��2�<q�Es ����kL;�6D��z��}7	ѩ�3�j3�z��zLo�[s�·B���Y��;:e��'���l�:Ƥǻ�#�i��B)1,,��(�2���k����=������Ž�n��-��T��jl���q�a����&lo;Ëo�0�GfT��V�h��:=35��>�KP	���P 7�K��kF9�{5A1�|���V(-C����7oa-潾�M�J�=S��K�Td�x���W�u�k�����Rw�����g��՘U�(,3r�'2Od	����1-qLf�A&�R�Fw!��Y�lse�
 $"nB�9�(�`�읃o7��@yU:<ʳ_�����	E �Cr�^��?Y��l�1d�)�# �� ���S�"rU���w�kن	�߃��$p�I�"��؊?��0����X�z��j<;���G�۵�Q���>��d#X�j��f���J\���N�u�=�{:�ޡ����.���=�}���nA7�qKV}-�2�'�C��W#�1�bY�z�8/��.	�:#���������p):F	��,�Qa�B�k%~�]w9�b_� *ք/*;#�X�*7������1V��NS%Zx�?�B��g���$�Y��6�1ſ����oO�e`s�؋�(��J5��S�M����.0X��E}j���s�E�_��Qx.N�;X�-oÂb�Ix���V���{�T��Zb'ͺ4]^��A��_Mz��L�*��b��"�e�;龯4%�JI�+>�(�/O)sa⼵� 3��Zm���;@l̂	2���coi�T7vj�#�\�o\��B�hm'��/�W�C����Mzڏ&p��#<9S~���#6A�֝���a%sVX|[d*W�\�� d[��Yd��Cy�3�����$�L����2tE�v���������w���)����;M�z�!�b��"��4/�'���EQ#b��\��Dnb��\�@+��:L��j������ocD��B��� �s2j?t΃3��Q�k���ȍ�����3���	y�w��7i1�42;Xb����\�3�A�����jf��[��\>��MP�*�́�f#o����ߐ���$�'�˳(K�y�춄��_%��uS;��[�ރ� .�VR��7�ׁ_T�7��h3��\ ��s9����斔�f(܊�STʼp���	�xK��
]��)�1�j��5u33�X&�.!MwN铪FyehXCDw^�$:1����{�p#��P�"�Zx�6v#>I��R�`�鼜�� <�V�jRrxQy�X�	�Z�����6�bG)鱘���٩	�@����%�,)��܏�����S!.�F^	w{qe����V�q��W-�D�9�8�2�=.�PQ�r��ݑ!N�����+
T���-��q'-�ÿ�O:����T��S<}x��P��f�F�:��n��g�p��u,����dn?��8�[_!�,Oj���H�Lˎ�G�i��j��!��C&�J��6�|�z��������r���zU�~(�Q$������ig1���Z�ScP;�Z���NҚs|9 %-���HV	d��Nq�M2&@�;A�2c~��w
Ws�ٚpuCz��MW�λ�ר1m ����.��Z��������h/����O�>m�5�V�)�|rQ��T26�;2c��4[�z=S�$���*��$s��V_�%�+%m�i�����4E����
E^�6*�Z{���$f�H�2��9Ml̩=k��a�LQ݇���}�ݑ}��Q.9:�