XlxV64EB    2e8b     cc0��:�܌�G���o��nf@@��Y��.7Y#�_S��9��!���+3��h�n^}�D��J`��T$}9.ȠV`�*F$�b�7S{��3�nXzڿ<�^�������T�i�B������{�5�`
(���������{V�G[+��>j0�뢹�^�N�qͣ\�҃~��u�.`޴b,�"�[�6塓����9��{_ݏE�~�y���͚��\�����z��;ߓD�= 0ى��`�Bm����{�7�/�h6N��N� �<߸�!�W�ٻde�0�#�������0�B���So�	��6�S\���X/lW'�Rc��ᄂ��*ߗ�q��/^���j2��1�q�yF]��=Ë�aϙI��o�'�S�2�����L�"n.��O�6�9-�����3c,��$��"�N��]m�f�R�<l�Mxqd����1�����;��YS���Q��~%7���Ec1K����I��$��;���4:f��ϴP3�� Z���߀?�D��8�����P�1����`��m@"�O�jZ���ڞ��äUp7��=g|e0���B��v��<ِ�V}��fm�~��z���rD,�+ֶ��g�9l�~�E��?+�?:�
�\�PU�S^F���Jnn��U�R��FU_��o���2��XZgOؙ��{�	
�d(W����&h�gn��ׄy��5.�OL����Y2�~y0�*�)c�:�	��jp0� �ø�@]�W�~���h�tvЖ �/�{����KJ�a�5]L!��s�>[��j���h��<i_�޹���I�u�J{ߥOs��HtZ���Y���:��QW�"f�j��Vaf��Gt�K�#��@^i;�J��7��:�k����!ʚ��D��������Z	�VuƵ�*�$���p��J�-��W�����p^�ji�
ȩF�c�4*�.���FsA>�E ���t޴w��n��2�Xbz���{�ӥ��>k��"�\�2Jd��j�4��DIG
�u�R���>�_��l�׀��8Y�[�M!ƭ���*����*In(ִ&f���"Uxㄙ]Z������.��y��b�6sD"���0_b��5�7�cH�deĺ �v���0�&BB5����1Cp"&?���+��^����gV�T�����J�uOn�	֙ޫH�S��1�	ݰ��\�E��d ǂ	m����<���<	�����=�_��	ӳ����Ưe�6�.9m�Ԉ�0���|��-�"qm�/��6`+i�ᴾ�j�"�"�e�~��*�\<Js2��=Pm*u�ۈxU]�}��!{3SM�R�+}ql���~Ѯ4�d�!��	;Mu�/�-���R�D���>ّs��^��`-cpЯ���w���t��IސPfx�u�u���ҵ6|_�3g�n���\�`ܕ`����l�&X������2b�Y�ÝY��iEޥ����	,�H���Q��ȭ_|+������Z�'�o1�\}s?��|�,��T�V��jwR�E[��@�N΄_�I0Kք��Q��2�z{t�H�~A]���7����[�Ȝ�� 5?w����6#瑻�:8�5Tx�m�_1�6I�[���]�|&烷��AV���������-�p���&~7x�6 ��	_�4|i =䐶����O�9Z�о���}��>N<h'�� ��O�6VC�- iv[�e�J��HW%������Nv�׃����/ɗ�V�Ud�ތ�����[�P-_',ʬ�vJiƢ�snz
�!pY]`��4 uTa�1"T_e�V8NXx��+��L!�@��V��z* ��!�r���4�Eε#R}e �,*�_6[	󮘕1��--�M�}��9��]`�A7�_G�D�ULA.kQ�R�uSG��-VL������뗙��ƉE�����He<@��&��置q=���T�Ɓ|�� ��h?��{'��38�
����@6�m��w��RtZ|N)�"��Ãt����Pu�!��W���Af�Q ��|m�'�cG{a�(P~�L~����N�`�5S�>���Ԋz�A4Syu��DG�F8�$Л;��c1����԰״O�5Y b��W�Q�ʞT�QQ{������׃PH���p})s fH���lGPC�V��������7����
^>~U��/��M�cY9V�g��c��-�=�񿈿w;|�I��V�Ց�gc�iI��1��'�f������â�U�3�8Q����l�\��d�1q}ur��>
j��.,Iኦu�B��ֽ�t��@;�e�eN��fJ�=�L9z}f��������`�	ʈ�� ��J ǒ�;����ge�/��0	p��Yt�,CFr2qFrG{H`��7���n�q30{�t�0������m;u�NX�����	Y=�e��B]��f�X*�xf�4!ߴ��k�J��@>����$�궻(����UC�BP[}ƳvQ�p@x�3`�[4;Z=�Ȯ7�SF�$��mT��7��ˡ�le�B�.ʧsxL�c���M��w*z���-Hk�H��J�ٕ���e�`�ZTO���p���v��3��T��}���_������>�5��Z��kh���lhLT��l`Nc������h�A�8t)�	)�n��|v��Բ�Ki�Y�k� ���p#�/�vx�z���*��$��R�ѝ�2�b�I5P���L_KB�³� �u ��b�����]_D�?i3׷��y�/�;�zsk�`���⍇8^�i`��r&(�L�+�r1+�7�%ˌ7���]�K�Ηr{��^���)gy� 9)�^Ch>oP�7��}MSA���u#�U��V�!ܿ�����߆o�/16��e����c�W���d��}{5��E�ʴ`�j�`M�2>� ����)�h���P�6LN ��tb9�8���trU��hD��a4��zo�%"�H�3�#:����&Ɉ�fI�w�<|�t��;VC����ߖ�j��Ӧ�� ��=?��k����̧8t���CǞkn����c%VE�ޝ�hmE�'�1�s�����X̩d!��JI7�;F�k��JS�g~�쎽�JDT\7���2����5q�g��%]�W�*J���A��_��.#L�tN�|;G�,�kp�^�H��窙aظ<�Y[gf���]R ���'3Ӏ�yIe��4�u�3�L�
���o�G	�ܽ[+���#l�LQ��