XlxV64EB    1ada     9e0�'�O��c�������7Sŉ��/�w8���'̏=dk#3��P$��4�����Q����i���B�C�'�Z
�6Yi�H	Rrl����N�i���1�_*L�e�Ld���x�Q/�kq"M3��;��c>=6�8&צ��o�bKOJɲ�1K2d��0�FV1hK�:�UM]@Ѿ���F.����w0C��!��8�z�]gu2�8�B���a���?A��U��1���}b����������R�����J��^�s;t�ك���p�b3��ɡι�YW������ȬFU���'t��#Շ�޵�>zX����8�k�ǧ�"�0�����6��IȂXS��韟�Ӏ�9���W?>��׏�${�F���VԱ�gn���V[��IU�A�%�~r{�c���H�U�����F�p� �Xs��
�ΩR:���8ҁ'X�o��jȒu��!f[��%rJJ��C"r�3q� iQ�t"����J�df,	��=���gү����b-���,��_�XbuSBu������۩1�p�wt�������!c��*�p��E��oOBegNDW�o���Z�鷤~yCk��	c��օ��ց���P�9]c����,w���'2���y���V��vN�/�����N��I&�đ���Q�^�>� n��L�ͫ`r���b߷H���L���z�gT^���F�\"��Xu������Q�y��2Ah2;�_�!OC�9DRc澰�!dP��"Ɏo`w���	���$��g�H���JsP��B��Fd�i�_�k�玴Uux:e1�>��(���ʴ��~:�/�ӈ��S,C�^��J\��b���ԇ������$`/��,&N�gO"���yE���n2��6��P��m�t������J�8�����(�{Xc��>4+$>e;Q��{Е�'7���&` N@���/�%|�:WOx�E����[� <���Y��A��~�����P	�RUT;������
:�1)`�O�t����kb�:h�HBL���v\[��G2x ��u����:�
��vb��L�r�:ȭ�R���'���:)�Cz.S-�q���
��[�Νnn��T����+���)�w ���LlS�a�օ�\x�*��ɐ;u!*;B��z�<I���Ù��vYH�<�נ��UA��D��z7�{��A��o��.c�:J+�>L���{iU�qI�~��2cRNǡ\f©-����1	�63k�Dw��^|�
���[���{��47;�	V�-�#���똧��M����YAk�)1�h�c~��V�z5�@b�$�j �'�~�}�G�����be�e=ƥ`����퉍����z;?��@�����w�R#����O��_"��yH�JA� �q��WP��*�-�l�l�zp�����Qx���=*��hf����0�DH�YRY�E.VD�����o�� �>Fp�b���0�í��PW�5-�	���Ʀ�����/*�)p��'��нN�q'���![�Q�)Up/ީCh*$i�B���b�57`gӐg��<� %,��1��+Ϣ�'ϥ�cUh%$H?�jq���2@}��䂠��-$��h��W��ؚ2q�R�n>Y��L�73�bt���Ec� ǧ<(۟EV��,:�;u�����:>8�03&�T���%��L`��w���i�Ѣ��݃ː>G.������d�sj�C�U���C����6e}�D�|����1�ؿd�`U7���]�K|�U��X|ڐ>qs�s1����}�`���7XC���{S�����O�ζ��1�S#y�m��[TT�fs�Y���?9/<}�jW�v�I������<���-��(.#�N�����p����mYd�C�N6� !H+�6>7������"D8Xɣ�ˇ�yi+-Ǯ��)��� ��W�Bj��ߍ�����Ua��]�q��w�`H�y"���)m���`���j��2�\ M�.��R5_��q��!�՛�p�C�cxO�<T}�����]�"6={Q@+p�,y-���0��Q,j�64!�T+�<K�x1)��_O�[�$��ֽ�!��Aױ�PH�cP��gVb!@�[�1��3�X��9I�G�!k�S8���e}J|���5G�\N����8a�Ǽ%}f��@\D������(����|N2�C�P�sq�h6��߉�L	��$�lE��[�C�V�թO�fd�G�5͐	^U�$��liI�/�@��_#C������ƻ��EC��F��kʤ�^�R�އ8󪊙�������T_����TT��q
0	6?qv�o Ԫd?�/�!���;�lê���(�FZL6~�o�TF��*�<�೬���3��x�#eCH���_x�W?���⯤�ʍr0��]T��=E�&�i\A�s5`CF�:�ŕ��>�V�]c��P?� 
ʢ�JW���G�v]���w�{�έ�2ݩ#r��1̱j