XlxV64EB    194f     9c0%����~�n�D�*��\̆�����-+O�b���n,ڶ�%�r�Gye�����>�s���X��4�3(�����G������c�m�J_����2)2TH�B°-&��g��f-�y�1Sڲ$̺�}�&'�nW1��c�W�!NC���s���B��9畛�����P��e�c�������������ށ�$����%�!A�ş�Ap���]�`=��c�ɕ�g+cK]��ʫ�~D@��?���Q��}0Z���=��mw�H!�/�+d�O��ʘ��,}��
@��v��z�'�tҎ�K�l����̞��0eÏ��^ �H~Y�lO]��9�h�(�ڜ����E�e��y�v�������NFv7$^R<�
�["A	�3�}7$�a��E�z&���يw����ֈ�՗_�'�D[�_�Y�&��a���Ms�G�g|�~�g�sP���k��n�M�Un �i(}e���&S�%.�0����-"���Le��o�����U��f�]3`�kp�z�����
-��qr��
��w�d�#�<A)~L�&pi�by�� ��k���x�ǺD$R&B
��E~	��~ט�K�m#�H0-�շK]���C㡥a�[�d�tE/g��w���e�(ʞ26��m�y��.0�~d7�����kX	�1~���|*�1���p���N��6�\հ�kb&�Lp'q��3���`�/�_��rHF
Ą��'�/U��e���>�T��^]�<�3���{ �a��b\�FN�1�e^�����\bU�#ϑȿ|:�����y���x|���%u��l[G-Qo�:ד4B��4��l,c�vG�Q�ًB9A����TJ�HM��Z\D��˶���֘��+�AD���Gv�eȧ��ӫ�B<'�����AUk$&�
�խ������n��Տ���ʪwEkƚ8҇��3#Џr=1�Փ�V��J�[rWW�Q��×g�Ȃ��W�b�.k�����i�g���]a��8z}1���������ɝ�B=��8+�~�����%T�m���h�V:�]�����V��!�[v�Q����8[������Za[9�0	=�-��QE$5�l)�F�~�R_���i�ĩ,�XSA)3��~�Q|�[G�f��}T.VX�/��k�f�@��R��cj���h����*����Vm��?^?ק] *>߈�%$��?��ϐ;�h�q���yM_ie1ݼ� �㋺C�����k��M�LJ���e�D��>m&��|��7�ء��&�¾���{%/�À�M���:����Ƌ�&S5	�9�,R���N70�?&�K�$����b����c��X���Ф��d����������S��-iN7�\��?����Tq��en�w�zRۇ��C7�MҘ1%;�@���1̛1�g�P�i��'v�n��(���oaᰕ�²7�k����Ӽ����M�\J̀����a�!��6Ǯs�V��IQ\k�J�3��˦��,ZӴW=��&-�]���<|�KK�o� �+R��qj �M&��Z�%�g�j[Yz��oSB�dh� M��_��#���֙�5ld���eQ������6�oQ-��/c��ܝ�T%��^W9}eZNr{{h|�����,�;����O]��Kq���=�
�|�p��Bv����0p�S�	٪�1J�4%iKMV�|�1��L�r�W���k&�Bhv�o�"����f���3Upes��o�n�����X4��FP�ɉz�7�����a�d��*�v洶�7^De��s@�l�7��#L�?��]����R�ƢF!;	o��K�JX���9��>�v�' �4J��uM���>U�G��5�s�A<N3�
��ì���Q?���G[���f�X��;"�����2�oʶ��d-�-8G����~��8��Dpǝ�"OU�t��L���ѯn����Q����	���ׅ���APQ��ȳ�ra�&�����-�7-���N^���ҸH�>�@m�|��T]�jb�����1����"%�L�J|�?���s����s��)��2v�J�_��g��|}<~9��/HxJ3�BEZ�2� m?Bʲj�a�̈́$�� t$��G�R�]7.����H�S��`�xZ���5�:b��O��JtD��H��|etR����܂/��?fq�7�N����#�3eS1}x���S�:��t0qrf4]U�	�ɉY�X��ʊW�]4�t�s�&{�w��o��yq�#���?����6����m����h����u�����ٰ��B�b�?ICV�jd���5�߉�{�D[������iw�#��訣�9�VK�r!Ģ~Qz���(�k�3/�a�z��b�^�)����
����6F�^�g�p=�m����nCR��&�'�vH��T6�KCp��3��0