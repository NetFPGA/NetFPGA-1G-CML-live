XlxV64EB    1554     7f0�jz�����7%�S~��N�?�4�Ij�c?��5�A>
ꯎ������������w�O0q��+R����O�ؽ�_t2��&[zXo��0�X��l���u�����V*e��}�T�NCi�����e�_ �f�?��%����&����L�|	/6N�'��rZC����V�� ��0����+�<T0�"˼�G1�\���ޠ����D�����0��j��|�����?>x%�@O�Y�nB�(\lٶ����X���<�r��`��� ��͏�����jޯ���v��:jA�9�%���zfP������(qe��A���(�&*��\�:0i�O�B�	?���w?��=��^�����l!��~E�ivL^��=�/Q!x�Y���Eaт��O�V?����&�.�o��yk$��v��^�N͹�1��o�$\��M��54횘0�ѓdD���5bh��o��ݍ�M�~r��J2�k�O��*���0�Q�>�]�"Z��I��NA�/`�(�NJ4�����̩(���]��ZUA��˂P�D��}�{ꆼi*\��	�?�5��xvF�<S�s��\�;Q �LL�eR�If.�O�#�-���zg_�#x<g�)B���Ă�ëwg�x���9BX���mߤ�.mq���MZ�Eqӹp<OD�U ��W�sR疯n��C�2��J��s�Tf�|W?�u�P��<�v�z\%��k)�b�����)Q?��{1��Y��f�h����)���F@����]��W��3ޖ/$��E:�[|����\�I����B�����6��'ֻ�P;��Wck z��ꀔ�������n8X�q��<��FD�P�~`�j�vlL��)� ^��t"=����U��!BͶ�B��|�2��ڷ�Oq�5)�$]��4��rl��������%U榁�goF�'�p��Y�EA6jr���^���[u�P+�9�%�E�Z>���[�SKwN�Q���2�
m��@N�Y��B�?�&���t��\}�xW~�{�2��7@nI��=ލ��C�x�i6f�y%|�5�4������2ly�+[wn
�Q���'əg���6,0_I�;��2��L%B�K�۾���,uo�� ��
��+�o`FՓ*��n��g0�����ok�d��-�a�	�ǖ79�{�%ͷ�R���_`�L:j��Q���ΐ��HiO�|��Kw�a`M;�1�>B��iH�77`��:���Xν�C�lE*2L�-h�G�O��sk}���ULe��h��C�e࿵a��X~#4+��ui֭c���o\"?C�F�&�����u+klj]��J��x����2����}܄�-l�����Yǯ����L;ڰ���gTz���ֲ�*0C����t��?`�6������]��}���k,m�OS�D[6Ð��:[q��7��p����k�S
3V����#���u�o!��d<���@�ʙ�itV�ph�4i��n�]���N,���{;ÄM���.�DXj�5�o>���_F�W���Кb�Z4���Ϻ���8��2~��%Gj���kڿ���$U��5��}�hu�F��a����Huܣ�j��0��Wa ��T<�ڻm$�@��)S�OK�.-�M_Rƹ^ a~��7L=PbU����л�4Y�}�G� *���L��1�$]��u��܂��&���r���ꊕ�]��i.��W���C"M
Ux�K�Y���ƭ_I���]n²�
ɛ���:<���L��"C��o�O3��{�Nc|T���ĒFIi)*�Xo�NG�z$m�2;N&�аO�s�m�"��O��, \B͞;��|��e�+�z��Cf�B��}W%�(��'%ఞ]��NڲO&r�D+�a{�?�sy��I�f$�,�	A"z�bˁB��3#M�u/Q��P�9˅����/����8	�}����,u�,Eh��ϝV��)5s�&@�.�u4��q�������a1ӡ