XlxV64EB    b718    1be0��5�!}C$�ʨ��
�Ql��j�P�՜��l�a� 0z}��\_�D@��}�kZ�Z1Ş�Jn�H
siY�5��Z�U��_Ɲe 9VNt�J�+T�(��h	-"����L��$S}{����;�?���rM�&����i�������?���5��;h7�	���o�u ���#��W��x�y���y������{pJ��pMj�qfG��3_�{:�P؀h��&6��+`>����9�~��K��'+ջ�Kc���g�w��:�Z0)��<�����)�)�]Wၦ��usy�����c�=�v
P��[w����mnk3���/1�a'��� �zi�7@����</��?����{�u}��\X���]2�UX��2��wm���r�#�IV�K��f���g2�Z�I��M�l�@O`��������4�ǆ&�,%�J]�}���ǅ��\�+-�;B���%SJ�L�r�[�]��l��q�+6`OC�#u�-?\�-��i/�C	�/P��������������������!��홤���QX�Fk��$ڝ�e�kde�҂x��/Rі������R�����м�	��^�Ox��C��Ι&��������sB�P_.��G�zJ�
Є)��ʯK�獹H����l���c�Oi4��gބ�	�);.r�,��U���s2Lз�C�^7U�5}r{�#�����Ƥ�H��/��}�>����>��µ�nw{���n��^��i�L=�M�O@�H\�s�Klw��Ҥ�o���]�Y��cf� J_�ę�=�O�+�
�;Z��tkW.�~�Ԍ�� ,��A1ޱ������{D*MOPF�t��,�񃹩F�)��4P�ګ0����!�t�F����O[Bԭ[������ G�(�m?���� 6i��9x;&y�5l�=t	�F�*�CJ�����3����$^$;74�Ԋ\��v��K�/Wg����=�Cd����*�C�V���(��"wdcS��^�� �<�#/t�q���) m�pt1���e�k�7"{v��
��ֲo��č�1J�-���qP�+3���W��A����O���YkYV�`�)�?a��C~DV�^nja���G�J�j�9̥��1� �}��������=]=����|�Ejx~�5�	�gU�ʷቾ^lp7iҀ}�;҃O?�~=��E# K��"FL�~���l<C�J(��A��mPr���{�C3����fm��tѡBN�f]u� #����?j����.�ȴZ%	��ݳF�Lt��M16����$���qbi��J%d�B�A��?:�3g`�.L뙲�dP�7j侶�^3Ml&��>���Wb�G����� ��t�gW�1��r���E)�A���J��B'������3FKs}�'(�;Wu<����0�D�J��֝ra)I��c�U�D�!��G^h�bx��d�z��6'�4���NF��ML%R�*t\�15\������?�6��N#'����7L����9LZ{�Z}`���W�]�'�$̯��f'�Xs$Rǟ�,��7ש�P�v�xތÂzV����k���Ә��d��6|u;j���]�)ސ��X���y�ǧ<!����7B�y(�+D�q扇g�5��n���ˢ�����)�*t�.F�)G�/�c=�NX��a�j���'��ErPck�sj�P�W�C��c�I�t���c;�>�t&D��g�Նݢ�&�}Ž�R�HU#xr�j�n��g�.������B{���-#uC�i�Z��(d3��)�T���Q'��/�n%��u��(0b�}�#$�V�Ϟ#�
�ن|A�m���%v���:�)���.7@��96Ep�^�b�ȥq�r��\8pj��1-����9wq���[e/��f���F���A/��7z]~�"4�P�ݭZ�q#�����I�	BB�'�����X�)9�ڼ	�l%mgd5����BR<BOvs6vQ!����#��ue�!)��ʧ���9��I�K~��H���q5$
p��La�c��	&`.۾7��ʒ�L���⡨���;2d���x�'��W���p*���WB
� �y�wC&^�٠j�-��l�o������'�ᛙ-�|3U��UƧU�J�0dH�����(���	P�_|-�W��j����9�,�>�<w� 2:.F����:��K+xzrݲ* ����m��Y�ֵ����?�	cA���֢uZ�����f�v��cq\Ev)�-��)) -S���϶���m{��������Z�8��"�!R��F@"Q���cXq&�ٓ��OM�<!8����
k�tOC��t=[;�b�2�h j�q�T���i�C���K��+��C��JFb������X�1��'�}�,����\�n9*-���*����X�y��5�k��AY�, y��ր%��je��iJv 7>��A�x� @Ҵ��W$Wgo`�r�3;�	�Wu%��[O̊X��dйe ����¹A|�.Qf�'���|�1R`��ԕ���O�Ĳ�:h^���˧&A�1����F�&����� 1G��DF���,�UL��JՋ(��lt��Wܲ�_qA?wu�������$xIۂKS��S6�x�ʬl�9=CO~�x{wk�!$@��qw�e���k�ߣ�,Jn���,-��������I�@��,�CE�F�h��3�������e\@A���bLXF����吃�yN.V�!��~��:������ѥV00b���������I���4���c��*H�vL��7�K��>�g˅�	7滉��;9�h�l��LLmiQ�ht;��*��=�I�r�8����8�iEL�>U�N5q�)5m����[c4�ξ��P-��k6\*��"�q�3b<�c>;.\�Y�`��u�DR���G��-�^y7�7m];!�1�h�#�"i!� Iz�_�|�8^��(����8�b?�j��2������ �p\2'U׬"��H�Ka_�Է�P��<^o�6v𘦢gq��!�	���#n7����H�����(��J�� n:{O�^�ޒB���U9���Wd�r�`D���O�'#y@�|���	���s���lZ�a�t�7��m����#V�.پ��*"��D��`��g�������en�~�!L1.;�@o��X^v���QL�ha?U0t����rZ�Y6�^`�f���x-cr@�+�("����si�0��X+��K�S�+��푒�qFF��_ş���]�#ε�ʬ�� ��Ȱ���H;o˛��ʃ��j���v"Lwk�+V69��8��-��'�r�c��.�r&�ϵ�)T� �q���V5`�\��DY�V�,��-�4$�ྐྵ�U̂}�a�%�?|Y����+�?�`=#����O�S#��e��k�u=/^�`��z��|v( 
}�Qp+��/���h2��"#����~�T*m�������Buh�r>��,�n���7郧���O-����_�����y���	�b�����d���-��E�ی��Դ�b�^�`���X�o�um����e�4h�z�����r�Ct��4x@R)�	��H�6��-s��\3,�Y���L^+��1O�� �}[��-�IL����[� ] ɂ�g;'�;Kί�i�#�zJ�ƺɻ���K(�rܻ��H�-*�")t�ǟ���˺d��s��8ntJ��h�e���*$�J��4�]6��,��0,P�3�N#�������������>��K�;>~ޡq#�\杰�d�a�CUgG?�Hk|;gR@Nۮ֒��8,8�&׬����b(��{K������(_�<��������él�����3|s��J[�&b���}K��(���N�MB��-�\3�I򤥛��c�{[��)Fa�!��u�.}�-1�hv��k�NjX)��	��50+�����U!�6_�&cFJ�~�y�bE��[�;�Ts�9�H}�B����7��mDL<ܚ5}�=�]B���9tZ!��:�l>��$��EU7��r��8�U+(9�}��26�Z�aȒ��v$|�Ig�I�w2z.�-��LH�+:�$a~�ƪ&L�,i_����FMH����@�s��<{�t�	�����р]�s���1�Fwz(���^^��Q��� FW�u!͓L�q4cS���lmJ�y;]�G���#�^�����HP�L1���SX��MY�-�(��̛�)7��b�C+�j��u�BD!�*�!���vD��A.�ێ?�M��S1���P5��^���~���J�kK.`�����mߢ~{��ه�����V	-jz�9K�4�
^��H���7�D�ᨴ��B+U��k�m�{�B���B�F��i|5�X',mt|fbך˕�E�Y�a�6���o���A�T�kfU�v�	}�a��r&O;�����~�?���w��r'��7��a�)aSO�����b����7������̘1����o��u���:<{��{�J=��������F�D&fJj�J�<;-ѹC�Q'7&���c�/K�_g�c��<P$�yP�<+c��D�U�@l����:��0_�HqP T��U��̴	m�ly�)��3���Xօ?_���;-��En}�c��������)��m��N1c󟵆�N��/*X.�:�.M��~�x�m��l��j�(8��\8� F��+��ލ���ɺ Iu�Y@�]�svx���6V�s�P���6��[�5U��ySE�wJ1r�e\fBN|	I�B���`�4g��QQ�j/���j)O@����3�𠿽�~nL��]��"�to����쑮@�4�L|�c�M�x�����IK+�ƱĆ[3�5���|�!��&����6<�q<����O�����vȗ��'2Ͻz�>���쩬9ȫ<��D5�e�7 �a!Z�y��N�~f��5'1���K�_l��OEHj����3Ff�l�`V�R�զ�3� Q7��c+��ae�X��+WWNf�*=~ �o;�4��`�)���M�p���ի����<����N�\4�	�e����-���~,�o��!J5�_��0[�;N��Z}��9F�q���x�l�����'�zV���1�3 Aw�-1��vR7����K��_�M}=����XO�g�U��'�4�S'1v�=@�u�ӬD��ݚ�r����xl'���h�72h@8g`5�Jr<�a��]U�pf�	�jf����ҙ��f�-����6x1��։/������%QK�;<�g�X)����1�G �.�H�G�d��ю��-P0%�qa_�(�,�2�]J�dJ�����5Lg�dN!ڞ��p�T��1���j�CSFE(k��!iD2������(=��`o'�����R���WD���J�Z:ś_V@`�R*o�,C�`�@*Y�k�������OW���<��a�9�7rT�dj�F^mP�u	o���6�H���U���[LXB� �L/Wo�u�(;"y9jl��u7j����/L���,�+�i	y-@�R Vk����R��o��gBFa��'�S��ߘ��X�%���{�h�s�t�����l�JX�<�j�A�X7�cx,�ɀ�v���{X,���۝g��c���5|@��Y������E��}-��5T���HKy#�6�B�����-�1p�R��5�K@���l4C!�kMe���f� ���L��B��6�9�����0�~\�\���GE<|�z0T����k��(aX���|��n�X/u�8ۃ��k#]��Ӕu�˫헙�KLz/��;�[�����ǜ��p�]�8r�>�
�у�
D�x腪���C��p1�&	ͦ����s5�e~�����(fSf͐!a+9N���2�0ׂ���ۭz��V+�G{�ke@��x|:��`�:,݋�P�ìҪb$���\xQ��c�S�E?	���"ǶP�h"	N�I�L�|�-e�:�@�2Cm~� �/�l�[���Y�cC�ao�������Uč}jJ^��0!N�L@Q|UКƸ����c��͟!�W'��F%Je
���Hhn��`��=p��e٣�7�ꕊ��� ����,-D���R!��Pi5S^������X�@-d1 F�[�s���~�s�4�舭���.N�Mn�P>�Q.pLqӵYRy� ����e�:
a�Ҩ��������]d�4uI�'{���� Cļ�+6�±��΋�ۜŉgt����ri���e��P�,2���A�Я�$ujT�G���y\B��J�$Ÿ� �:'+XG�c�Ӷ�4�������~!<8
(�Irј�9�@;z�;��ۭ^��]�,�5��T�CYr~�k�Y��y/_�D��aW/r�>�~��X�\�-�vc]����+���-����rp�C�4?�!����)����60F��I	����n�ni�Xd���U`牆(3:�(�g�v��誚���Ъ��s[@�:��	n/1�<�~��
�mA2����;����I�t�/��W���,&�$�>Kk(��\+�mg��&)��R�k�b�g0f��1���UR��V�H��JE�U�P������ճ��6�Jk�V7|ԃ-w�zU"�f!`JΟj2[�	�U���1&�k�TF�p1nmИ��9bt�]�PB���ƲvO�Q��J;�0*�3d5�lgu)ƝK$)�\]�K�$�J^�&<_d�0��8X�ĵ�Ftm�r�
����+Vh���{-_.a���_1�Ak�1�x�,��#C��cm9��Yoj��<����}��M�d��s��a�
l���_�y�Uǯ��#�)j�`a��Nd�,0���#���EC�Q���/,��)���9<,�;��������է9ø�oe	}C͔Q&���s��RsDLW�� �A���7���sL����r�����'��x+��4��Ʌ0�쿔���2de\