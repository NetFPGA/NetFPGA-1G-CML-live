XlxV64EB    7282    1750�l,����oA�	H��3�V�jdR���8P��q
�K�L�����,�G�'�� �/"�0*��F�|�:��8}�V4"8S�3<��J���ԏ���T]��;$�`��*wG��X��Քנy��M�uw����d��v�=t��%k��W
��?��+�x|�}-�2��*�L��&�V�i��"v1 %!O3�Ĕpm�z���XMj���%�bH�"R���E���3���fX(2R ��������$���HO�)k(��JQ�g�2ڎ�s!���2��9-N����W*J21Jؾ�"zcv�S���u��9���5�|�D�pϹ	oq)m���n�y����hᇪ1�Z�c�t�nK��}�+�F����J׶��`ᠯ4_��Ws:����ʬf�l"؍^LK��܃'�s8�,C��9~vS��*C�J�B.A��������sE��l-*`���(���I˝�|��o,}X�/���~�ԁ 2.�䧭~劖2�W����.������#�\�-���Fł	���"z>k�H�{-\0�5��O� l?|L�5Y���UE��2�Y���#�=u�	_���iz�L2lI�.D��c�X57�O��V��4t�7�2_�fiw��Z��H�`�	ZC��C���EX tI`��J��x�c��C�S46��m��?#����|�2T:��zc��Z�g&j<����:E�3(��̾)7u��4=| Ȏ��0Dd�:��C
����=~��}����>����R��p�VK��j{?Ks�*� �>Frs�T�`���ٱ�-��_���%�ҿ8䋪��YF��B�%Z�<�,���z�R�����va��&7I[��%]��XM��ݻ��`K@������]��� t���N�2:����Z�S@f�{�}�zP�f}�4
��˨Q�y{�ᨩ8�QUƏt����<i��qtLt]݅f�Q��
G����R��i����z@ڲ�w��Lɩv��08��0�{$�6(�r��Bk�+�Ŏ����3��g��pK�
6�b�C�&�5�ۼ���8sB�5����]B���E���x/Q������h�Z���w��!E��*���ґ��{G���Z��>?�jz�t'4S#�x�n�_��p�A�\�+��Gox��$/K���{]��EZ��$���0��]��OZHV����G'V�I�LF>����qIݢ.3�u��z��[_�uNB�.mR&2vX��K���J��7OZ��`?��y�S3}:�ᾂ�eե�L��^��܈�ips|,ṹ�/�NU_v�R������{�t\��L��Q�a�$7 Gܽ=�?�����"�c��|����[�����!ʥ�/W��PG�m��ؗ�sX��;���ePH�(�5g�&�^٫�c4�h|v�������ot�{x���K���[�뾅_0����'<�Fmb��APU�ЬD��!
�� vկ�/q�+��^��#��F
���Dm��v��ː����1�HVg�	�w��=��h8��(Q��g���(�կ/ �����՜��n܂���v�]o��Hϲ��*�C|9Rm6n���%�ݨ�c�HV�P�S��"
@m'V�1D�n�0�����9����wȖю �ϖ�x~��w��3q����oF@�kF��T.KJ�����^g�?	�����s��-F���'��e��)r�l�\m�VXȝ�w�p;�q�$N6�Ø�ڋ���u7���<���?t�^�H�_.�>?2B �b�"O�U�?�8d�%r7E�|�aS�sTl��$M��A����kR 95k���z�����=��K@�O/>��w,_��T�mn?��H����荚�x�0�Oߊ�J�;xӃ���a�@( M ��4b�e�Ib7�sM�|���G3�5b�����@)�6���H������i�3��E;P���+���z�r�������i�oy"}^��J��B�"�[Ѫ�u���y(��MI�i覘�"%�8@�`�n`U�щ̖X���!���`�
�Q�?���FabE~cqx1*�E���`�|�Ձ��� 
Z�|�X���L���r,+����F
)��;�sN$�y��69��-�)�'V",U%�~����n���X2��W�����:gK�_M�Ca:G��M �v��Zx����-o�L塋�,GZ[��Gu�W�W�ۈ��T��-�@��գc����?��4&�p���	l�9͔$�@7����A�$���5?@�lL�ͱ�1��mi(�]�tC���/غ�p���yV
�Ň�N���_ѷo���%n��8)L1���}
,����`;L�Ht:�:O�בK�H��k���S8�~{�di�&0�i9C�?�I­� ���;�#�2vLy�H�4��3�[�e�OI��xY>	�Ŕv�+y�(2�-�<ha�Z)s($2X�rG���?�ؔ�8�.֢ܼ���9�����a6�����Hy.�/�P��\$u3���i˚��p�XU� �A|ltI*�1�ؙ���t�H�S�wޣ^��I�Ư�2ʸ�@��$Ο<�d�k�wm#EjU�c�I�����e>X���4�[�9��VV	~yN�pi}$��֥�(� �=f��-�M&x;
)���Y��v�|���3���Ԍs\ݰ����}g�ۻ����t�Yc��"���_��A|r*�\m;���j�SuD��r6y��AC��(+#D�F��'����O��ܺ3�u���I�6������Wb���$"c�ୖU�}0�Ⱥk�0t�6!v�5��W��C�b�ϙ�b2��7K�e����C&O�*� ��q���ѱ�{��g~����,������.�QY�1�hj���p���!̂9dKF�R�m��aw�#sS���Ͳ)�˳�O8�T�έ�M��x��nm�}v�(Z,�����f�����sP����_<�<��4�a�L��d�ԕ���Y��ZO��$
J�)�~�r�Xؓw.���:����gW�3��?�5��Ƙ(L��}�e����$��(Z��(��Aŵ#��X)�G��j��:w������j�3�T���a�o"����0����C�0�2#��(�.`r���,�#�r�h��q��}�1�`��w�-%����~��\��#�fy� :�(�R^Hu�*lL�C<D��CL�z�P�]VnA.Mԕ������A�
�i�8�+~h޳x�O,�Q��H�9�W�.*�t7���Sx��A�siBq/?�����J�]G�B��;j)�^d��U�����4l|�Y��QI+�O���wv���H�W�!9������s̘BP�u�d"�cr"%��[�x��x	�k�q9 )��J;���N�y����HRi�?3�ĂΩ��|"���vڤIq1l�(�Y?9�@f���v$�P�c+��<-��wSR���{E��+�t���ap�����Z�`�߷�v�?"�A%�k��K�3�(�Q��f�/~��tam�L�8o8�j�2��:��jdu{����!p���K���`���D�j�.�R:D�ZqAn&�eȬ6t �J�4c���Sy��s��|p�ؤ�mL��1g�@~�a��� s@���>w������`�I5��4|�E��+��Nr�5У^#-��Ⱦh'r"�R�j����^�_�$�a>�R)���f5��/��J��-�1cIPԋ���
��@�V��J�W���L;�sn� ���t�^�!d,
�f�+��͗#O#ZY���K=U��{'|
�Lc�,Z���^d��}/�����Rd�lU�8�"vv��w�j��=>�c��u�N��j�����.���Trᚚ�G7�1����wA@�����ꂴ*�U���51�w@/a�H�PDG,�i e��ֈ���§�­��q�*�Ӛ �ק>F_QP��t
)����t�?.�Ռ,L#BK�R$h׿"u������+������3Z��_�{��]&�^�&v�Q��{d�o3y�6��.W��Ԫ���g(�ĔA	�a�Q�l�Y������S4X�|��88���,�0*V��DôRP����"(�ߔt,v��@*o��r��d�e�,���$���='"��G�!62_el�d��Θ/�e݃���l�v�]?��l�G�Anb�0�4es4��.��J�$�Bh��"�K>����'$��{�T#^�,KZ�����; TN/��lrq�{����H��d�5�to}t���C����]s�CY���l�ל�����V��9��븕��@���2�͒7��[��QE��D�i����Փg�w�
;=����g�`��n�G��j�XcT��o��2Y���A�&HC�u�F�Y`�_~h��zדs��S���"�_���iP"����O6@m�O����c�ab��D�R�V͙�,��K6"1s6�#�}�,
����H��znt%#���\lf*�i�a��y��ƞ:p�L�4����vA,���b���3"�UF���ly�Lں=���H�.!��nqg����z��;y2��D+Y/ N�8�)-P¾�r��Y�k���dz���ΥL}bP
��T�P�T��he����V���t�F��|Y���ݳ.�D;��/���?Q�˗�^�$������ԃ��j��(�x� e�jǿ3&;�>�����_�9$�ˇH�mc���\�3��BW
�tR@�ӄ�.u��v���X;Q	�˻�ɧ.ݥ�C'�X4��Ui�6c@���\�94��E,���4s<h�8FJs�<q�ӎ���������`�i\���#k�3����� �� 7	��_r/�6]y��n�Y�&�f���ڐdS+�hn�Np�6S؎����H���-�[x��7���(UX��с���]�ʘ��bR8�a��IuЁ.U0s��8��j���!+���y�vP!���;]Cv5�h����c{�F��֞nB ��ϱ���t�e���۫W���b�_%�q�beEb!�@�]�]D�D�5�k/F��#����P�/P�غ<f���x|�H���X��g �֗�
��� �#��1�n�r��|�����_e��8�Р�Lb:�ݮ�3m�r>�G��G�asp��@֫����*���ƴ�_����_k�M��v��)Y�O�& �P�Q��i%���:�D�Z��,0#h� �`���_ �Č�l���H��)�\�,�'HSNl��!��[ �&��۩`�e�B��G.�b�7S�0{��z�%�e{]=��=7�9���`��z��~�2?���OP����*�ZA�i��:�MJ�f��fl���D�ٜ\��5�a��J��;�.~��
¬]��F$�K)��U<������������U������Se{T �Kl�[NK{d��Q]�i�����4�*a9e�:V���@������Sc�y�b/Y���՚q����6�"��K$2{*�]D�Ql���`U����l�KI���,��ڿ ٬�D��V��Jz�o�Xζޭһ&i����(B6�D���n��[[C�l1����H����L��E� SR��r�_��O����$�Ng�����Pޓv
X|�����1ov�c96O��Y� ��?��mA�R��ӒW2h��y���i���U�9֕�Po�s��9���_mr�'O�ډJ�[��.ܢ�.��x�a8��8V�ղH1���wڔ�S@�.����l�,��T��r�4©.�zfT�٨(5l������īY/�4 �K!��X݅������Ԙ��)�4���Y�`����X�I	&}ʼ�׸ʎ������UdQ��^��5yR�