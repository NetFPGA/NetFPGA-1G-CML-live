XlxV64EB    1648     880x���]-@M+*̔[�r�5<q�q�I}�p����C*�G�.EGw�o^ݟ����_����n۹1!J���w_k\~���BN|N������V7]�b���6�C�P�6W56S���,N��o��^K����|���ǿ��j��։̏�k�g�ђ]���n�7�����U�w��s2xP�:,�h��c�b8��K�T�����QǬZ�0=������|n��f���{>�;,�i��1/��20�/����%�7�Z0d��u��%�M���5��J%?��&�9R��{�>F"j��J�J�6�&���������(͡��?����!�K��ǬPJ"�R�/V[�K�=9g�d�|�`����_�U�"�F�oCj*��D8n!Kr�j[��{���r
��)^]�uy`���������c%����m�&/�I�}*�����ܱ��e�k��4�0R^��m�:������:�2�1zۧ�a%ר�� �H�B�������Lx�R-+cy�����ܿ�!����,�����U%��/���Ɏ4{���+��Ybv�������O���ߊ��Ŵ4}�[�#�qAE%�din���DY�T8w��'ߓ7ȓ	;oF����p���\����.��å�l��SKg�2R�≞�
���ϴ�f~amSK��W�N��{�9��V�̍h)WZRI��*��Sw��ݗ�:i��z1/�Q/��6�}�xB��E�v� �pӫ�prQ���g�nq
Ȓ��E�\vxNFv�N�j�&Ea�d��a܏+V������g��%��=�?��<Ub]\�����P���)z��|Z:�
�c�o��������6r7KV&U��a����a�J�g0m�����2�r���%��.���a<O���V:�<^ɢ�[�蘁@��`Dq~��<���� �׮�,x�~*K/�K�b4�|BjT�@�2�z��Lg�^?_;�
U�O9��G��~cz��4RE}�?0�@fhL��9����,��<g�É�~ьqDO_��Bs;��_?�me����5��#ѷ�7 �sww�F��,�81�C�"�{r����̱۠�ZI[�.���C�>�S���?�C���@����$�"]	{J`�	�2m��Dt)�(R��6���Yg�D��B�����9��dݖ8(]���}X����9^�TJ�vi"+ꥤ�ݜ;�I�	p{�
���L��g�˹~���yB�e�'��6Wu������/1�]�%S��<wsD'?uJ��XE���k���P�sq�]�<S#�vr *���;n��VO�VKi"Z���=����W�m�	�����Ex�5�����{R0e��#�_y�F���K-�ClL�Ú�[q��t�h�&��Z�z�Xb�wS�:"���#qxA#y��@�m����T��bo^I7=:;P�� 5٬�G�ƫ@��K��f��c�PP6�̧��*&�_#���tH��}"��X~�Z���2-e���6��1&�,��/�4J
�u��,��-�fܚ�&鿖���R�����!wh���I���𠣛)${`1k�JH�5?���Q�H�9vA�I�mq�ބvĚ��Z�l☘�>mkF ���Ӭ��W��oH|�UQw�恁�1VQ˳b&5h�۩��:�� ����C��J�^<KC�����q�0��\;�5�x6��%o�/���c��&�3�ł������V@u��@��<T�	w���>*f�^���x��C��O����UDc�
�^84�
��D��5��Ȁ6�#~"o@"��^����Rhk.A�k��S��_O0e���� 7bxbg�4g9ю0Y�{>(S�����A�qL�m�+��߯���5�q��z����f�W�);��y1�\su�u��u��e��D�s٦��G� S�x�Y�j�G>a�/��>b�q�'7�QL9�?�ln|�a�*��(�uY7e�m½c�\��`Qu�5����~�'��������^���d�ޔ���՗vi�X��$�� �ܞ�묎��_��<TB��� �V�%MW�Q0�R��R�����P���c�-F�����O����xS�\	K�j�