XlxV64EB    1f78     9e0�a��6��aJ��T��	z3PI��֑1À��2R;�t�Z�n�r�'�;����U�yL�{�M@Z#i�x�E�8v7A��RT�42Y!��I&eՓ�
>�G��M�y�7ѽ��{�Y`q:lL��?p��̭�#���5b�>@��F#Z9+{�n�ε�&��JH�f��ֽ���a��1����Ɇ$�F���-�+E�Nw�U�����ީ����a�_Њr_�8��k2ʣ�|��J������f��`#��]oL̇�����b"�W���[�湽8��40x��`�ܟ���=B�Uw�����\��{b,--�H��_�ب� ��G̗b��J�4F�QT�п5RJ����h�?o��N7�akϫ_�2��˩����Yɕ��>�d��i�{ӇEnY(z闓��L!�Nrfr,�n�k�����sI�KH������!}@msg�d}sИr�r����X/`#wDP,�wy�ڞt�;IP���J`K�nFei����#s�	0�ܳXS�Pfk����5i�N��8lW�$��c�s�cв.���7մS��>��6qVgk�S҇NZ�����j�Y�h�з>��s/<`�b_,zħ�זP�	���l�`���w��#����~}G��+S��s����m��w�'�*(We�|�j�Or^��C���:�=�8�	�b�̱\�ήѝ���͹��T�t�J�.�b�����f[΅��x�F�<��:�%h�T��*����uZ���LLsX```*xj2�%	bD�O�#MX��}�#��)fU}<f��<�=�k|!T�|�tU�L,��A�1Su�^U���$���R;�����Erh���r; ���C~�u@XvS�r ��~o���������Ʌ�LQ7=;�hhL���@` `z�o��&M��v��[X�:ڋh���.r�
�KG[j, ���I��&J�T�Wk��T8^^�{�}Z5ڰJa����牡����[�AS�a#�GP$�Ʊ������
�Ya����d3��}���t�»�6F�R2�CS�D^�4"�����$�A��޸�jk��D���P�.b��ApU-��"�ˀ��(��/A+���F,K�J ��i��&"�s���tu�d}������~�ڗ�
�W]T
b�;	����Aj��N]y��iܜY��轧�h)ܸX��U,^���c7�֓FK�,��;�����0�\n��K���}b�L{���~�.�$���ͻ���8�lG;��C����?'�;��619k��U�O�l:`�eQ�ϯ[�0�H���K�fk��r(�:/��2�_��/*_����,�<Wp),C���!���iu<qO��������K�y���*b-+P�R�! GH�	݅�-�PT!�B��X�;�-�EŹj0eV�'�2�&�	��sT��Č���g�_=9���Ԥ1p�	�j؟���[+7�0)uf	�޷r3�x�QSQ��O�Z��o�Cԣn�b[JaY�����9�fA���P-�d�jmn�j�S��F���a�7��%^j�\*�Rv��''
 �`M&�_
d�\%tyUS�t8�<w��Ũ9��$D1�)�(�.~��Q����
���U�fĳ|1~�P3��E�x2���KVD��¡��ە�]�ً�S�Q��y�����ZY��E���D�90=p��!��؝�6CS��,eڑP�<�=J�-��N�@��Ƞ\��J��)5�t>$h�i	���蒜#�>	Y~���84��GO�Ȼ��oq�v�G�f��Ēy���c�nd}�.��X'j�����{�wF���k�D�^v��H
�Y���9��~:�+���OPV1&��$ʮ-���=�_s�1�+6���.CX���83���D1��1x�'��4�&�q�c�}䒽�4>��u��J�eP%���REx��h��IY��p�Yq��]�����:F5�.`�T�C-3�ĺ5>� �I����Dr^��=�Ӛ����X�TkJ@0S��zz��Qo�GdI�7x�_ْM�n� ����y��ԞbfU�~��ޅ�%9�)K��s����f�Y2��-�}��f��'�?��pv�-
�"V� �vu+p��|l�L��0gϷdy���Đ^�~m7Ǝҽ���j%x�g@���M�}�Gu�[�T���e:,є�L�9��LMeبk6��H`]q���&�J����O��HS��+�),O�4a#z�������)Qoa���Q��9}��V��G)�V����nTѽ�8̶h�X2R�Z���`҃m�pH���ġ���b�s�M4S�u�G�KɄ�c�)��ը�њ�E#���;���b�AUf����"���O���dJn�/&ۻ8��V�f��TV�&qY��m��l�7��X�q<��}R|���3�?Ϲ�f�< L������*DZm,�C/��'�A� z�����p�$�w���$l�u�no���