XlxV64EB    3f9b    10f0-CԼU�x�(� ��U(�@�4)]���sg�GֶŠ����I
-2bv�E�oZV��ZN����4���SN�a�pI�6�^뛟|�q�L@�2�C��hc&��gTn�?E[.�f���0Ңݵyp�C(��6A����t��+ԀrY-�;ٻ
�������#v��ȿg�^ d�'��|]�Dӫ4ۃ�SmV�
�
E�xZ3�S)�Q�Y[/�����~��J�+Nv��Ͷ�E�_�!_���'i���pd6��"�N<�|�\�{��dWV!D@|�f�C�.<���!y,���V3����\�m$e�L�@�CO<�$.U�^��\[''���9�MX�ʍyM]m�&�(�^��8��+��`$WV�$^X�p��u^`�M�*k/B�����)̵m��<H��`H���'��od��6�'Nm��C@xb���P��=X�K���;����?R+"���-l��3�l�OH��iR��Hm��Lސ#�*me=p������Q���;�\-�.nM4�brcSLRċ���ƹDڐt��
c�)���2ٕ��9�(?K�!��1F�#7�4o�wS��+����_|jM-j2oR��G�r�#g��m��3�S^^)pG�c�H<�\9g�P���﫪<�����qa|����3�kx��j�1��4nZ&�Q8�u�t�\8�[q�0_D|L0��\ ���Ň+�~����-' �!1�Xķ\'�W��$��v/P���'F��`���ìR�1�z��G��zʻ��2M;M��C~�u��lZ��\oiz�:~��H���כ)�9��������\�Éa���NXbK;���11�7o(+/;?��ҐZ�?�O_]_ٽ�[��7K��ſ�&W{U�
L�Mo���M2�tz�y�ː�4��?�O�Ѷ|�Kto	Ң�@<��VR#?� ϊ��:�1I�l�y�I(�.���T�%�Q�l��Q=X=^����*kc&If05O0��뵱@��N�
��H�e����P����@�RAlL�E�Ϳ�'n�Q)v`�%�?)���СD�CR�Ť$i�bEIDg{�^@빠7��~1�t-�v����b?�z�\�(HJ�~C�NY3��o�ڄ�&�i[�S�ն���i���.2!+�oV�Ԉ%N� �rnZ��p{���)����S����nyѯ��i���E	��h$a���ED#�&�{�sx�7qh��F���l����n�e��e/��~�vow�־o���Nu?��W\!��jt��,MƩ��V�5\]�U>H�W7���X�	�s��TF��M���
����%�糑�^�x��9�	�i�鹣Y	�,>� J����ExoT�?��B��T,C�b0F&�۠�]3�L��[7�U�=d��iˍ�v�=%�P�CVkd�4R;�����?E�67��1@�-Tj�E����l�j�-Uq���
<����Wƺ~�U+�D�֭�0=�*��Q.���4��Ru�L�I7&C��_B�d���]qrlo���]׳���=օ���;qA�_��`����[��@���kbǎ�%��M�p�p���^m�,x=�Q�Uv���a3t��@+K8.�v�%�tV��T�J������M9��Pӥ2CBM#��y�Z!��j�͜Q{т^���\P���f�/F����I63����?(@��,�;d���A��-V�A�P�I
OB�C2����T�-;Zt'��֐�X��A+��!���G�}��5egK%C0�N���Yi�0#0O>N�e�~ �M#�����n^s�d.�Mf$ ��U��O�����	�L&������Z2�:l�R�4W�� ��9_�赢�l>�&5@�]�Y8�oDh>�,8\u��vAf��zbf��&lo��xv�N��9�xC	\e�._�m��رᄡ
�\���U�J�w4�<�H�����
�fDmA�J����nE�,むF6��fX���tSml���%�������O����s���$�\�#e��~/2��a0�K���I�'�����U����IK�	a���E�m�ʑA�v[�)ֈ�e�е�xV�rj�?9]qr �*�(�4���=�ݲ7�^X��Xl�E<�K��8?�>�&e3�KuH?v{9�e�
�Q�ċk���N��@X6r�\����n{�AM�e���~n�����w�M�C��n�<���<�_�#"MN���C�A^Q718��^;��l����6��5��T�\F�q3��	3�td�[�/����t|���{.^�mL,�'��� v�ve݀�Ё�y����'���U,֟
f����2��~T}/f�J��L�����5D�y�*G{�o^
���3��4ǎp��<��/�b�ze�E�����~���|�Y�������C�Q"V��l��1p�6	�Y$��#m�P�m�@^Xm��!���tHx����S
q�h���"p������˴$���W��+��\
¥�10���K~��\�e��ir�J�-7)���()aл��u�e��F�d<[9P%��mQ���$�o�0D��=+�I�9�"Ty��7�&�ݤ�\����`�>H�*?�{Udw��ϊ�/�����qr~7��qg�F���v7v��@���Y-��ώ=��N�p�k�Q�6�7�Fh�".3�ϙ	j�vf��9�,�5��' ��e�������ʩ�#�mR��ZT���O�'uпrx~1qJ����{  ���0�3w6�~��)SJ���\��gQ���y��J���M�q )pX{��]��$!"�����ִ�ȬF����f�dl�0���
,sH����pvpmф,��j{�> ��{��"�S�� \;���wqO���ʿm�g�^dK��4�5�p�N:��$5����19�o�팣����v8��M��'������߱LI�c���k�Pɢ�9'�l4�>^7��2,a�d�՟�|>ǌ\�ς	�ꑁ|��͹��쬴�04i�3蜣�R�3 P���o}���n�&m��� 5��S�������;_pNX���bV���#h��Ou:�@gԎ���[��K�͹�=�U�\��!1�ZJ�$Z�/d�p�Yu��&��n��ȁ��͎�y����ȕ��r @�(�w|ݛ�<�A����5��1$Cљ���x�@d��h濤��h	���]6�~!d�����u�k|jղ��*w��ˠu5}��Uv��c�pl��G=mo���Ӿ�������1�*p�+iO�VN-���v�3� ��w�o�����i�0M�,˅��d�y�dG�œWV$}W�|�QH!���Jo�Ȅ���^�.��~7�?���G����r��li�Q�������և�Ʈ��&`��u�v�5Fު���}��yS����G��>=��_{�<FT�α� 7�և���ð2q��/m+d���Vg��&���y~]�d��h����?�#K���C�����~õ(�����!pw�ďbA�_ ��{�k����1�0�6�f�I��K�A�8��%�t7P�腐=�qx��@t�;�_��H-%;׻�ٌ�÷�W��������S�5��E�m!�M�Va\Kfpg%���|P7l����޺�)�9ˍ�����X��F�VRCxC?7�јMi���\��+�.8R���c�/�n�ì�"�ZY����惥�g ��"	!Q�ou��l�`����g���������(9���q�kt��lD9șռHЗr�=φ?�糍�$��� yv�{e7u��:�[�a���}��	-�?J����ݦ��wƭ6�����C�~5��h߂w4���t�9�M�P?��^5r���/K]�D�%��֞TDb��z`"�V*G�2�?�N��{�?⻯�"D J>80�Ϙ觰���V'�@0��G�+���x.,�ܦ�%�g�485�h�x3��Q�ЉT���s9�ڞ�O����h��12.(]��|��+�v�R?�υ�Ճ-)��S�|��>
)?�G��tq*��$+>z��a����C�1R�l��i8�TXv� ���%��l5�y/Wg�bP�A4�b.O[<w����**Ojrs��a��*ܫU�%B��Q����o��U�9�p�q����z��@�����4�Hh�4�����%Ǌ��e̔'���v�L�zw9�Hj��߲��+�����Ӫ1�A�%����j���5T���(	zd����e���\���{�:z�Kd�������D��I�:��