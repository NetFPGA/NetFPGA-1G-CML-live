XlxV64EB    3b27     f00�Wf�B
��հ����� ���h.�
�z�mbK�ڧ��nC�c�8��4��p������2�{�e���o]��(��0��ʾ�x��D-��n�waM�Z��}�iJ:A�`W�'H�ξ�S�y��e��0��Q��W�V솆6ɘN�9�WL���&K�N���	�Ë8e�|��RߓXh8
�c��(�����W ߃�NG@톸��p� [��I�1��l��H�D��߼��8�C����=�U���'��s+�����z���&?b�H[mG��'����-�\�(������]0؏]Ǵ�LNC)Fŧ1�@m${�����ޕ��_����[I�O�SX��z�����x�?
�,�d�n؞���d^�e�B��_�]Ïm3�ᯎ�0�F	�C���1��+��?����\a��"a+Y*(��zj����?������u
�� `�x����1!�T����Y������cz'��PN� ����)?T��e`��E#M}�mm��ǃxCO���)ײ��{��7�$��#�b[���t pX5to�(g�����q�x�����_��O�k[����)J�)6�K����=��7��FX/Q&z�gV��!^/�^�� �Ե��<��p� c����d�0����;s��*��ܭ��ڣ֑�|"��0Z+_c�C�?Gh���=&,�f�yu���D �)�J|J��ϩq��3�^0��p��c�&��o[�З�垨�X�1OO\�H����C T�XN�U�_���yK\b�%�;�z0�ᖞC�;S0�hYxX�.}���@�L�84��}4��Y`ؙG'Ƙe�+�(���r��	�y��aW���t�h��U@ñp�-�4��:�J��zo�3L�yi��޷�?\�h��.�Hq����Ó1v���|h,��7v�u�n�O��E%��a~���`�B�R6T⹐�ŧ$�ڞr�wn���O�R���h\�V텠�5*� �������_cuϓ�:��E���r�A�x=�P�<r/BO�=:��
Ѓ]z�"U��9�SF�!+u]��&!�2��&�s'̡����᱂�j����#e�\^�+hkv�c.}1b�(�W�i���+�%�IY4��;�x�5`�,>�{S�~	�&{�#Ȯ�4�S{I����^�mP��A�������^��@ ����Y^{�	h��X����J{��{��z���6JC�|߳1�	r���v
R#8+R�N�0Y� ������鋚qG��4�P1^������tt�X`�C�B�^-���� ���ӳ�4�= xI�W�מ>�pJۄ�ʽ�Ӿ��#�+@7�]ݡwl���8��3=D'��V}$�~�,F	:��B�U������R�>�t��NH"D�믫^=^��rIe�f�����/�STN��AC_���[M���	��|X��.�|ӊ����Rw��Ql/�aс�H|��������K���4X-��!�"�u�wo,ؽv���z+�]��r�k]�D]T(ą
R1P���Y؃}��C+����m��n����ܦ�c#�����{(}�Ȑ�d���qWP�@<F���g$[��~���f�p��Z���5k'���*[�X���_qloY��W���|�rv�����}�6�FF�n����� j�D���z�n��a\螘��՜pC�����l�l�x�+�_%�A�ο��E��5^�ŷb���2VL�$���0��4�����L̕	Nb&m3�A7�9���/�d�i�J�̂m�W��<y�����2�+B�(qu&�P���@Ȕ�N�z�'�I!e@	���@V;	AOd|(��h�ͧ�I�H	��Z��|W�ݷ.El�}�:���8k�`����5ָ��bC0����j�����L��d9����x뷉��	t�K�i�u��s��vs�)��f���91���!����~W�%�|0�a꿔�k[P��ڔ�kb�
�&���SuQ�|^���ͷ�B�l���a+ݧdp�@j�����5�nq\���L, 本p��L8�E�Zg���yn�h�d����m �=Wd(����:�r�������{C!д^�9���[� �c�Q�)��z:�#e��ٖ�|�6�a;������-�������J���g�}���ص��T(9�m���9m]أ	b�"n���tH�q�p?]���	��Uc(-�?&PjR��|���e�&{	�_��>����=���[Nނ_�?�Y>����7�p�Q�J�D�5�N��M��b�S�x4[}F�7F,S��Iq��A��������#ʋ}�֔�М��k�T�N�ϴ���^*�$�z�X���)�u��(�oףKl!yJ��|��&𘵟һ�Ai��#�0[-{���V���2��[5}!��N+EޔT�p���=ȅݭ 1�W�Ltp�&A�0KaKa�#cZ�ki�*����H쫦�U��+w*:XȈ��f�0=~P�]}�EO�t��n7R��ܾ�g
����Y����&[~�5����3'4C5�xݍ�쉗�'��]ʐM�>��ޚ�X�oQ&�O{����J�L�U�2 ����2�n���Xj��@'h���R��z���JH��8+ܓ�Q��P��*���p~�0%�yS} ���c�`-���)�Y�[phh3C/s}��_�ة!�Z�M�����&��F�����{=7�5�֙t�[)h��e�P>0}�D����&�\�o��;;��̙�4EFE"Y�j��mT^eTm�m�L�Z��>���:u�Qx"35i�/�(bvы3��c�EF^��YҨ���C�$�9�^̓C��	�F�,G�Qձ�qu��DϚ2�(�%���U�>�m�_%E����(�����T4���)���P�����sw2<n��׬1�nKNd�w���B#����(=�@���[<D�d$[�@ZU3�\W���?�;M��R]l���\������ƭr�����쨎���\����uF?��&�`��0���*T�o\@p�=ݷ<z�k�`9�.I�OW�\�odH�~�r`���d�kG�֝e�wa�İ3H�z�H:�#����J�i!�M'��C��,j�1�FY>/�ȟ�)(y�oԔ,矫����t��MLS���
�h�3����@���_�o��U�H8�$�R��eШ���^��Lk���R�˂�	�6��$z,�w֭��+tA�&�f�dt��K�� [N�ץ�mR�M9n���B��\�9T�+9$F����<2=����D|���i	u���8*uX�]�mh܎c�[ }�Z͸ǣIl��MtO�OO����Q:!�Q;I?S�$���#�M/�*.�����>=k��5���J����g�Dűu��xh�v�31�Եn��n��RN�E�Ŧ<[���_(Ǯ:�R�fE���͝�}�	�yW2�����s
6��J�-l�'6'���yN���_���-�1jXDx�,�ۯi��8h:ؑS�~^L�]�i�bR1J�Lz@�R(�Pss�X�>�P��kŅ�NV����B^b3�`6r|���a��g���B-����G/�]�ߣ���h5�,��;�9u���ǜT��*2 �B��p����$�1&����UJ4��Tl�R�NM�;an�0^�O7ī�K�(����1�d�Ԓ�q��E��zZk�پT��,Z�{RCT/<Cl���VR�u�+ٰ�r��q-I�o���v�h���n�d��a��1}%L