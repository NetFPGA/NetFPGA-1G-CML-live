XlxV64EB    28d6     be0���4�A�� � �Ͷ&Gޅ��tZTҺ��L�z�9����H�AI�т?����UK&��+����wy��V��rK�Dv��(�Zs������閁����d�dz����{>�V֨E�����E�$�V��꼤�a�����]ς̣?a({��X�.���Ԡ�-?��}��!}�t�����)X�Ι���Ϸ����Ɉ�mj��rY���J�0���>~,"g �����~�ze-��q[�ҽ����Z���u����c5�\����(�G�y�"͑yy�h>M ���r<�G?W-�G�j���E�7 �5���C�G��	�[^ �;Xb���1�߇��N@�����aJ�E"M؝-���۪'x��<w�����vf�U^mDq��/3��p���#�܀A�y7��?ǂ�q"�辳)M���ץ��q�n�h�kg�>ṪJ��.4q� � h���a�Px��E�·=Ϯ3Hd����l�H�Q�{� b�eɓj�P5��Ҁ��se0���w��۔�Nal������`�0�����,X�G��J:�f���a�Z��¹1��EK���)R�.\�u|5��i6��1YD�8�Rq�bfZbzu��%�\�7	��xC:��^���2`�^:I\����b�Up�SV��rJ6��$wG�U#�X��}G���ݭ�����Fe/yMYK�bHW��@����K����]D��&k�R�}�	�7�7$?rq����/�Bid���� [[y��scB�"A��k%���Qmc@�4N��{���7Y؟��Q)W �2t��n��W��3��Ĭ�	hV�-�\��*�4~�QLz� ��5�ʲ�j�̞�VwW�O�~����b6(�pa��>���|����h��n��ж#э��\|H��w�������wNR�Z֬R���EU�h��	���|3[�5���o����}$6<��m������1��cx��6�q�c����-�S9��$jBb	�;�0!'܆1�y�YN��EO���7�$Ս�O�V���V<󷲁�c'��I�m8�?YWA�`zQ��ѠMt�Z١c�>�0�P��ldR�`��=���Ν������x�g�|&۽w��yTk�#��Ɵ\`���j&|���ѳ��|����֢J�y������aw�-��%.��s��+H���ݟo�
�.�pwO)�x���;��W���O��k�Vl�ǻ�J�57b��RU�����iZ��N8�؂;��/�H�긚[k��K#�
��K�k�3_oN�n.��M54��B��< �3��9�6��
�7]/��Ќ���u��5�a`	�0Ƚ-1�F��>Rh���������n��ʮ�k��S�0Z���*�bWX����^�+�2����H�q㕨�$�Z��\��&+�k� �^W� 8Ugx&��o��c?�?6��<g���,K,��o1�>^��R�
�s�Lxf��Fb��ٰ�g_8^���6H�Gb�Ѻ�_��J�M�`�����]��^�#�|�/��+�\�#�W����Qp�ZR���lF<�Րy^��^�'�����98��\a n����{!`s��:<��T�s��X/��g��\[�L��1��������u8Hi&v{@Li+�N��u�e���M���Ɔ�Ӏ�X��J��l��ԾH������Y�{k<w9�d��Q�����⌦���0�]gUx�1O&*Y\��+K\�9~Pڇ��*F���t�!����, �.S��c&�*��(�J:��� ��kq4��9�1�5hǏ/�+*{&�W�d��eeH���1a�j�H#~�وp��H`:��3t\��η!ȗC-@ׄ���������%�Zq�18��{��rRc��o��d�㕵� H1+a����
�/�3��y|���e���n�K���,�F����=\6v���yM�oz����(���#��r�� �Q�����΀3#���T��Qv�D��b�QZf�ٹ�O4����P�ɥ�.?�)`��/�z���R	9���v����x�A�2V��N�z*:�2���CG*�֫�uG�hsR�0R�V8�}Ya�K��r�%��+ؕ لԔ��]�I�&B�K�O�F�Y�k��	:>�"�܃��O����F��8:e-f�2�x�T��"����>3ΞP����sƔ/E!��<ާ��C)Kx,:L0�,8��J�+e'����.T��V��c5!�������aP�/��u��x4���l�ϋ<�a�f�G��8����S�3����-�/vjo]1"1iV��Rݤ�x6e��ux��������%Qc䓥�j��悽����Df���(#u�@��8Hx�S�h��� �Ff=���+7���B	���'��
��T  %w��	m�mi��ጢl��p��g��p"�iXc��U�{�#�����u����3Z-<�%��z�A\\�$X��ǩ��gR+�R��@����R�U���BU��&W���t�xlsc����G�{�1�w�3Z�����J��H�����,U+ӹ�����L���%pS�[,���Oȴ�y˗2*K�z� H��=bc�3��RؾFe[qlX(x�8��,'n��d̎[+�������;�ernnx�6���J3�T}�۞����=�I���˨����pk^aN�#���$����ļ.=e� �1b�H��4�S��uS��	�[Fa�>5�`o�q��S��U��e��z.��Qm�����>���*�Y����9͛k�'YY#kq�x�݋�	�ۛ���Wl�^>����4؂�)�]S$�&O�^䅭�1H�x���)i��{��������UߘSg�_!yN�~Zs�"�ts1��M)Q��VR��X����|蚸���M��vVD�,��&w$�f
�)��#��^q����n@��4��\�=i���;�5����_���h�kU���L��