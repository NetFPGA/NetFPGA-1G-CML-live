XlxV64EB    1d2a     9f0h�V湼�~��q��He�|�n�w����hD���~�z��;� ��\��T{1�2ݏ|�c����1�����lI�lQ{��۹X�o��w��a��o�ɜ�91}�- ��F��+�� �X�+�7;�b��
�4S�{A{�o���i��ާs�I��ǀ�I��g�����`?SM�U�C����ze1�4�Ϡ������
�����K`��/�oq��1�"3�9�va:_��G,�I&��w�~��2�-@�ӦP���-�(��s::k��7��R3�ņ����;[C�k�竦�(��7���h�n�ZCDZ���d���TU't�5dm�:9x��<Fj�3Aj�d����i ��۰�}�I-�i�l��� ��R�$#�@51[q�V�Cj*Dďo���ru_0kP�fǦ��v��wi����ȚK�~n>~p0��_o���_n��
?
o��*�Ev�w�|h��B��.׳l.�Q����n��\�@MAc.���	 ���P���1�h
�cs�i��g����؎A��ڟK�9���A��q�{������N��f\���xAb̪�mF%סPf��̋��%Q7I؇<��1��VYm2S��N ���������6��|
�q.����{�3/c����8�SmH��8��̥2�����:v\�^ypis`�:I�����m��
1�^&aV$��
vPC� RϻRӑP�����T�Ι�ʷ.�V��|�l##�� �㴶�O��ޖ��gq�����
�#SYd��w������$-�,��3�mtT����Y0�W�k\!ؼ����0�����Q��X/�n��*9��߹sߐ!R҉�x�
,�*�i2$��o��΁��'�8�5z�}�t�	b>�"�p���6.Р�o i/�ST��+k
aN�:#sa��]����{��5��9�*:O� <E���C�^�bԲ8�$J��jJ���J�~�����9F�q/���w^�Y$,�4�RV���`e��O�"��H��Ė��E<�}�Iڐv�M������w�.�KD�#�Á\�����rz���5$���� �E�m�E���r�S�hy�
v�y�4V�I��YM]hK}o��yű��� �8;;٬��fd��3��D��	u��;��\8q-�J��/!\�3�Kl�nV�9[gVi���t��(�/�U�]J�u$�
e�!j�;ʩM�*Q�(k�3J�~��	��{��%��:L���ˑ���	����5�i(��s�\�*2_K.��6 ��4]2���FH�_�0����<'"�3�2�O�ΐ�H;�
��+��P/�������"K�;���$Bk��j��:@�g�v�E�͠� ���D�r)V�b�� -�_��BW�P�pU��fz��$�������*�-�K���Ԕ���m|����Hgͭ�R�D�����ǚ	�U�dɸ№]����l�b >1����0(攍�o����}(W�R-��?Y����+7d�8(�QtNo������f#ϮZ~<Ϫ��nDy����kP@8����(�wPO?r`���p94���%.G����Z����(Y���4���>���O�+��	hυ�3�
;�Tu�g��)�
%7�(X��9��3��so�L�d��y�y��+����­��UY��Y�W�aG�΋�@��H�
�堍i���RN��u�$��7��@�5��I��D�jg0��J�߻;�ҏ"C�3�6;�q&,��U&��h����������\w٧U
��yIF�����tQz�g��[�"$-���z�X�f'���T���[�
�OO1~��⋢��a�3˘%%.�#�:�� .t�,N�i_r�L�v9n؎�6XsѠ]6!<��q'7�/�Pp��	i��P h�7�>�gi���ӯ$�CP?B���V�v�q����9L��L5�\����q���&���<���T"���?<t���i%+u��@s�B*��p������0��_1�>�B��q�Uۀ�ͧ�e,�"ޫ̖����?��z�>��j�q��M�Xs+�φ��M���W�5��9��i?��K���]q��6c!�J�*p���$I55�(Q�N���ZL��1�E��/<����EW���bқu�����-���Q�L"�Γ�ҒX�L��*3��#�|���KMb������n�q9�S�/ܩR��-'r��
�A��1���J�Ј�^}/d��C����ѫ�	�s$���� �a�[gWֲ�m�����jP��g/���6[�|�&s�#M�_0�M����Or9���lax�jnި��TY�������j��s�A��'���'�[?�uVf� U�����1V@[)VQ2<@��4���S/��҈�c�C�Y��y�J��.� �R�f�6�@����*n��,���pH%/��~��Fl�87�+±�h��Ov-�X����5��@��)c��