XlxV64EB    3f2a     fd0 ����Z}����n�͋mk#KÒb(tf�^*P��,7\_d�v��@9@����c��G��o�*��J93<�#J�O��o���D	�:!�ʯ��|�ר619�4���/�j�Q����&�S����&�Z��L��=S6fIx��w�oD����@��R��*���q�5������X�+$$��Pyq���=^��y;s��
;�iF��N�Ûk�t���O�WyiU��ΰ_jɎn��J�wO;4؊j�E�vI}�@�� ���u���=�7 �(�5�N}n���
��'�#r����N�'3	񲖉�gQ�	���R,�/��V�v�&�3z nc �0���d̃���Kj� `��i��*���@�-[���Je�c�.n�-�R���|��M$��ad�Ɂ�Z��* 1��R�+HF�x�e��{���W�b�Z��͋�/�Ϝ8�9����/��%�M��8�＝��x�;7ߞ�R8@g!3�mi:!�7&���@�n�[����v�Y�'�����������j�ɇ��Z��}���*��[ig���Yy�.8O�7s�\����*�P#���!��Rf�є���2��Ŀ>m��ʜ0{��V�}�Z��^�S!1�%�ߜ���j��q
F-�΋�#[o�4��a�4)�E=	��o��
vh�h��m��C.S�K�[�J��j�.�/�JțVޡ)�4uy��UW�G=�����Y�h�y��\B���(����CG�3䬣��;� �ᘻM[��ڪ��r���&o=_����߱��Q��<G`�3��*D��GR}Oc��U�(vku��Z���A���G�T�V'���Y���aA�2^τ�s�Q0"q�z���u�⽯V�6�M꒼�w�cNR�6�ё�]v�x���_��{�e��&�GU18�D���gՑ�l�M�o� X�K�����\�ӵ��܄l�p�}�t�q��2,��eO��n�Ab���"U��J��Oᖵ��$¬���az��NS�d��7�+O��Ւ<7hUGJ�������'OW�z�"<"�[���
��ݳ�{�
�C�N�����M�� �И�>)��*�Mðne��G��yW�<�A)#b 9�#3f��ճ��(j#�k2=�M�룋���e޾����qxL)�9�X�Y�20h�[���j]Zq�h1�vɞ_Q5Λ��e�&49� {�Co����{�s17�T/�X��ф������O��e�d2ex»Y7;&�B�̋��|��h=9-d��P���ce=��+�mhN�VP*�!>�A���\*mؤ������ﲪI�7���!���W��0x)��:$�N���c��1�������]�6���=�? {<φ9
�(�8�c�FzK �N�ze�\!~ ��v�Y�}q<ċtH���=b�*����Ǥ�O�^�����TѢ�c�f(���XFM=��g	���c#��?S�� ���f�pV��D�ۥ�dr��;�B�z�Wx�<���<�K$��[������6�S�v.�$�K�QaV>~c��$���I��p���4���v;	�!��̝�@U��|qPH� ���?�W=��j��K]�3��ǎ��C&g{\��'�RL��i�T��㞻��h��{9����m%�4���>��R�<4ϋ��7`�⬊yf�Bg���@�~�
{n�A+��7DX��n��=�G�)���j�G"p� Z#SJM6]W��-�I�ɨ�8,��ւ$@9�!�Gò�E��z9�.���q+�Τ5#bݘ���V_�u�<S������>�*k�>���j��4�L��O��:{����I�9�Ϳ�ԢqF�tD#��ْ$�c����n^��W����u��-�V�!Q��[��~:�'LR��\z�]T��<* Fi6
�/%���rG!ιU*��~H�j��݄�k���/��w�4u���"��\�4�V���X+~	K]�@��"<o<�T��:��j�|$Ȧ���;���%i;�����:cl�X"F������FI��#K [b-Z&�<����Q�iS�����
4WGT���)�~�իה���G�j�6L���cbX@�Z���Y6u�&�������$�3�}�S_q~0x�-���0g̻`I��~�%�b9����[V���K�1�_�ZcJ�,��L'/�۩Np�K��l����I�f��L�%�y`D1��˩�+	���M#ia+'r��,����u��UL��X3�\ʢW��||�?��}A��^گG���]�Pz�I���a&��2$���|��e����#2WD^�9CY�P��0�4	�s���r�wB{~���U�:��?�9 �����&d���(��5�1TB�Y$�JH&�S���b�S�b�]�W��O�Bc��:*)�^�bkφ(I�i.��D�1Ln�����?SZb�5ӱԼ�T�i|5�2oZ������*�a��*���+�~�1���M9,x�Y���#�_��N�l�_��#l�{�`3\h�;�ƛ�7�-S�-y�l���-�d"-����>݋=`̜���w�eRwV��`(�5������A7��[{8I.��@[$7����gw�^���>�Ĩ���tC-C�{��3���H�PW ���G��!��%�b,�����N�'�V)M	�;C��+�p��s��X\����g�W&����p0���!���G5�b�e�r��-�C`��Z�E	Y7��֥�w��p��Gv���0[PQ�?��\h4-��%���j�1��T�L]O[(�j�lt��j«�\&
��u��N���dK1�o����tZj["t@Lh>rb�����C�/;t�}3خ ®>JE����=B5ٚ���'�`�xe���E I�t�x�gx;�~�^Rg�EK���U7S"g���a��1�q�Jt�A���Y,RJ��,-�}C������<KM��9,�)fi�-Ux���4c7��1��A�Fo�<��:�
V3�v���Q�[>w�^�u)\�B��	�KI�zn��|Vp6$cr2L[���œv�[�'c�Փ��/0_�I6���W�KJ69W�BO'�Y��+��i��,��9u�����Vfu��Bƌ�g�"��>��"���}���A�N�L��=�r��b[2�$I�W�67EH���������$(���R�E��%��Ԁ�i����I-���p��2t���M���\�=�ť��vOQ.�h�����0*������4m�-`��U�
��H]���&�*B��A����)%fz����:&�"���J���"���iW	>ߔ�QԸ�f����ǌf�~8��(	��7�+�F��ި!3
&��>k��4����#�UM������Y�U��n�0�u��n5Q"I��S�R��X�6!�d���;(��l�:$*4��e�zuDD�X���d�:4,R��d����
��~�a�5#���8ȷuCl|I�k��f�G�/8J tN1W���k��3~9�Y;]�w��Z��B!��3u��c�T2L*LI�q��'�C����:}GQ�)!v�".I�E��#:�����Zp�������W�ǯ��E��s�jHn�Z����z"��.��]Z�
'�qۑe�'O���&.��ٺ�T�+Ȕ����U��pA���i�t��m�|t:��u'P����,f�e6�#Bq@ !kz�(�^\�Q)ؔܣ����3J���n�S���^X�����������Y���d�n�Jƀ^
V){Ep@y@��s�<���\��Q���]DGThu p��Ȕk-�Lle��l[��(���U���QrJ���䆧)!�a���H��-����j���)5X�o	g�8o^c�T���^�(#6�����U�{O�+ʊ����
��a�e�G�0�dv�����{�j�g˭����m"�q�z,����ј^1t�▦O	�2͖���;u���>L�-? �2χd�)�