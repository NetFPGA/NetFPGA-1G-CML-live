-- ******************************************************************************
 -- *  Design:
 -- *        NetFlow_Simple_10G_Bram
 -- *  
 -- *  NetFPGA-10G http://www.netfpga.org
 -- *
 -- *  File:
 -- *        hash_function.vhd
 -- *
 -- *  Pcore:
 -- *        netflow_cache
 -- *
 -- *  Authors:
 -- *        Marco Forconesi, Gustavo Sutter, Sergio Lopez-Buedo
 -- *
 -- *  Description:
 -- *        A simple hash function to allocate the active flows on the flow-table.
 -- *        It is made using polynomial division.
-- ******************************************************************************


library ieee;
use ieee.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;
use ieee.numeric_std.all;

entity hash_function is
generic (  
  INPUT_WIDTH : natural := 104;
  OUTPUT_WIDTH: natural := 12
  );
port (
  hash_input  : in std_logic_vector(INPUT_WIDTH-1 downto 0);      
  hash_output : out std_logic_vector(OUTPUT_WIDTH-1 downto 0)       
  );

end hash_function;


architecture hash_function_arch of hash_function is

begin
  
--autogenerated
------------------------------------------------------------------
-- Conditional hash functions generates. Depends on the hash_output width
------------------------------------------------------------------
hash_funct_12bits: if(OUTPUT_WIDTH = 12) generate
	hash_output(0) <= hash_input(0) xor hash_input(1) xor hash_input(2) xor hash_input(3) xor hash_input(4) xor hash_input(5) xor hash_input(6) xor hash_input(7) xor hash_input(8) xor hash_input(11) xor hash_input(12) xor hash_input(13) xor hash_input(14) xor hash_input(15) xor hash_input(16) xor hash_input(17) xor hash_input(22) xor hash_input(23) xor hash_input(24) xor hash_input(25) xor hash_input(26) xor hash_input(29) xor hash_input(30) xor hash_input(33) xor hash_input(34) xor hash_input(35) xor hash_input(44) xor hash_input(47) xor hash_input(48) xor hash_input(49) xor hash_input(50) xor hash_input(51) xor hash_input(52) xor hash_input(54) xor hash_input(58) xor hash_input(59) xor hash_input(60) xor hash_input(61) xor hash_input(63) xor hash_input(64) xor hash_input(66) xor hash_input(69) xor hash_input(70) xor hash_input(72) xor hash_input(75) xor hash_input(76) xor hash_input(81) xor hash_input(82) xor hash_input(88) xor hash_input(89) xor hash_input(94) xor hash_input(95) xor hash_input(96) xor hash_input(101) xor hash_input(102) ; 
	hash_output(1) <= hash_input(0) xor hash_input(9) xor hash_input(11) xor hash_input(18) xor hash_input(22) xor hash_input(27) xor hash_input(29) xor hash_input(31) xor hash_input(33) xor hash_input(36) xor hash_input(44) xor hash_input(45) xor hash_input(47) xor hash_input(53) xor hash_input(54) xor hash_input(55) xor hash_input(58) xor hash_input(62) xor hash_input(63) xor hash_input(65) xor hash_input(66) xor hash_input(67) xor hash_input(69) xor hash_input(71) xor hash_input(72) xor hash_input(73) xor hash_input(75) xor hash_input(77) xor hash_input(81) xor hash_input(83) xor hash_input(88) xor hash_input(90) xor hash_input(94) xor hash_input(97) xor hash_input(101) xor hash_input(103) ; 
	hash_output(2) <= hash_input(0) xor hash_input(2) xor hash_input(3) xor hash_input(4) xor hash_input(5) xor hash_input(6) xor hash_input(7) xor hash_input(8) xor hash_input(10) xor hash_input(11) xor hash_input(13) xor hash_input(14) xor hash_input(15) xor hash_input(16) xor hash_input(17) xor hash_input(19) xor hash_input(22) xor hash_input(24) xor hash_input(25) xor hash_input(26) xor hash_input(28) xor hash_input(29) xor hash_input(32) xor hash_input(33) xor hash_input(35) xor hash_input(37) xor hash_input(44) xor hash_input(45) xor hash_input(46) xor hash_input(47) xor hash_input(49) xor hash_input(50) xor hash_input(51) xor hash_input(52) xor hash_input(55) xor hash_input(56) xor hash_input(58) xor hash_input(60) xor hash_input(61) xor hash_input(67) xor hash_input(68) xor hash_input(69) xor hash_input(73) xor hash_input(74) xor hash_input(75) xor hash_input(78) xor hash_input(81) xor hash_input(84) xor hash_input(88) xor hash_input(91) xor hash_input(94) xor hash_input(96) xor hash_input(98) xor hash_input(101) ; 
	hash_output(3) <= hash_input(0) xor hash_input(2) xor hash_input(9) xor hash_input(13) xor hash_input(18) xor hash_input(20) xor hash_input(22) xor hash_input(24) xor hash_input(27) xor hash_input(35) xor hash_input(36) xor hash_input(38) xor hash_input(44) xor hash_input(45) xor hash_input(46) xor hash_input(49) xor hash_input(53) xor hash_input(54) xor hash_input(56) xor hash_input(57) xor hash_input(58) xor hash_input(60) xor hash_input(62) xor hash_input(63) xor hash_input(64) xor hash_input(66) xor hash_input(68) xor hash_input(72) xor hash_input(74) xor hash_input(79) xor hash_input(81) xor hash_input(85) xor hash_input(88) xor hash_input(92) xor hash_input(94) xor hash_input(96) xor hash_input(97) xor hash_input(99) xor hash_input(101) ; 
	hash_output(4) <= hash_input(1) xor hash_input(3) xor hash_input(10) xor hash_input(14) xor hash_input(19) xor hash_input(21) xor hash_input(23) xor hash_input(25) xor hash_input(28) xor hash_input(36) xor hash_input(37) xor hash_input(39) xor hash_input(45) xor hash_input(46) xor hash_input(47) xor hash_input(50) xor hash_input(54) xor hash_input(55) xor hash_input(57) xor hash_input(58) xor hash_input(59) xor hash_input(61) xor hash_input(63) xor hash_input(64) xor hash_input(65) xor hash_input(67) xor hash_input(69) xor hash_input(73) xor hash_input(75) xor hash_input(80) xor hash_input(82) xor hash_input(86) xor hash_input(89) xor hash_input(93) xor hash_input(95) xor hash_input(97) xor hash_input(98) xor hash_input(100) xor hash_input(102) ; 
	hash_output(5) <= hash_input(2) xor hash_input(4) xor hash_input(11) xor hash_input(15) xor hash_input(20) xor hash_input(22) xor hash_input(24) xor hash_input(26) xor hash_input(29) xor hash_input(37) xor hash_input(38) xor hash_input(40) xor hash_input(46) xor hash_input(47) xor hash_input(48) xor hash_input(51) xor hash_input(55) xor hash_input(56) xor hash_input(58) xor hash_input(59) xor hash_input(60) xor hash_input(62) xor hash_input(64) xor hash_input(65) xor hash_input(66) xor hash_input(68) xor hash_input(70) xor hash_input(74) xor hash_input(76) xor hash_input(81) xor hash_input(83) xor hash_input(87) xor hash_input(90) xor hash_input(94) xor hash_input(96) xor hash_input(98) xor hash_input(99) xor hash_input(101) xor hash_input(103) ; 
	hash_output(6) <= hash_input(3) xor hash_input(5) xor hash_input(12) xor hash_input(16) xor hash_input(21) xor hash_input(23) xor hash_input(25) xor hash_input(27) xor hash_input(30) xor hash_input(38) xor hash_input(39) xor hash_input(41) xor hash_input(47) xor hash_input(48) xor hash_input(49) xor hash_input(52) xor hash_input(56) xor hash_input(57) xor hash_input(59) xor hash_input(60) xor hash_input(61) xor hash_input(63) xor hash_input(65) xor hash_input(66) xor hash_input(67) xor hash_input(69) xor hash_input(71) xor hash_input(75) xor hash_input(77) xor hash_input(82) xor hash_input(84) xor hash_input(88) xor hash_input(91) xor hash_input(95) xor hash_input(97) xor hash_input(99) xor hash_input(100) xor hash_input(102) ; 
	hash_output(7) <= hash_input(4) xor hash_input(6) xor hash_input(13) xor hash_input(17) xor hash_input(22) xor hash_input(24) xor hash_input(26) xor hash_input(28) xor hash_input(31) xor hash_input(39) xor hash_input(40) xor hash_input(42) xor hash_input(48) xor hash_input(49) xor hash_input(50) xor hash_input(53) xor hash_input(57) xor hash_input(58) xor hash_input(60) xor hash_input(61) xor hash_input(62) xor hash_input(64) xor hash_input(66) xor hash_input(67) xor hash_input(68) xor hash_input(70) xor hash_input(72) xor hash_input(76) xor hash_input(78) xor hash_input(83) xor hash_input(85) xor hash_input(89) xor hash_input(92) xor hash_input(96) xor hash_input(98) xor hash_input(100) xor hash_input(101) xor hash_input(103) ; 
	hash_output(8) <= hash_input(5) xor hash_input(7) xor hash_input(14) xor hash_input(18) xor hash_input(23) xor hash_input(25) xor hash_input(27) xor hash_input(29) xor hash_input(32) xor hash_input(40) xor hash_input(41) xor hash_input(43) xor hash_input(49) xor hash_input(50) xor hash_input(51) xor hash_input(54) xor hash_input(58) xor hash_input(59) xor hash_input(61) xor hash_input(62) xor hash_input(63) xor hash_input(65) xor hash_input(67) xor hash_input(68) xor hash_input(69) xor hash_input(71) xor hash_input(73) xor hash_input(77) xor hash_input(79) xor hash_input(84) xor hash_input(86) xor hash_input(90) xor hash_input(93) xor hash_input(97) xor hash_input(99) xor hash_input(101) xor hash_input(102) ; 
	hash_output(9) <= hash_input(6) xor hash_input(8) xor hash_input(15) xor hash_input(19) xor hash_input(24) xor hash_input(26) xor hash_input(28) xor hash_input(30) xor hash_input(33) xor hash_input(41) xor hash_input(42) xor hash_input(44) xor hash_input(50) xor hash_input(51) xor hash_input(52) xor hash_input(55) xor hash_input(59) xor hash_input(60) xor hash_input(62) xor hash_input(63) xor hash_input(64) xor hash_input(66) xor hash_input(68) xor hash_input(69) xor hash_input(70) xor hash_input(72) xor hash_input(74) xor hash_input(78) xor hash_input(80) xor hash_input(85) xor hash_input(87) xor hash_input(91) xor hash_input(94) xor hash_input(98) xor hash_input(100) xor hash_input(102) xor hash_input(103) ; 
	hash_output(10) <= hash_input(7) xor hash_input(9) xor hash_input(16) xor hash_input(20) xor hash_input(25) xor hash_input(27) xor hash_input(29) xor hash_input(31) xor hash_input(34) xor hash_input(42) xor hash_input(43) xor hash_input(45) xor hash_input(51) xor hash_input(52) xor hash_input(53) xor hash_input(56) xor hash_input(60) xor hash_input(61) xor hash_input(63) xor hash_input(64) xor hash_input(65) xor hash_input(67) xor hash_input(69) xor hash_input(70) xor hash_input(71) xor hash_input(73) xor hash_input(75) xor hash_input(79) xor hash_input(81) xor hash_input(86) xor hash_input(88) xor hash_input(92) xor hash_input(95) xor hash_input(99) xor hash_input(101) xor hash_input(103) ; 
	hash_output(11) <= hash_input(0) xor hash_input(1) xor hash_input(2) xor hash_input(3) xor hash_input(4) xor hash_input(5) xor hash_input(6) xor hash_input(7) xor hash_input(10) xor hash_input(11) xor hash_input(12) xor hash_input(13) xor hash_input(14) xor hash_input(15) xor hash_input(16) xor hash_input(21) xor hash_input(22) xor hash_input(23) xor hash_input(24) xor hash_input(25) xor hash_input(28) xor hash_input(29) xor hash_input(32) xor hash_input(33) xor hash_input(34) xor hash_input(43) xor hash_input(46) xor hash_input(47) xor hash_input(48) xor hash_input(49) xor hash_input(50) xor hash_input(51) xor hash_input(53) xor hash_input(57) xor hash_input(58) xor hash_input(59) xor hash_input(60) xor hash_input(62) xor hash_input(63) xor hash_input(65) xor hash_input(68) xor hash_input(69) xor hash_input(71) xor hash_input(74) xor hash_input(75) xor hash_input(80) xor hash_input(81) xor hash_input(87) xor hash_input(88) xor hash_input(93) xor hash_input(94) xor hash_input(95) xor hash_input(100) xor hash_input(101) ; 
end generate;
	
hash_funct_11bits: if(OUTPUT_WIDTH = 11) generate
	hash_output(0) <= hash_input(0) xor hash_input(2) xor hash_input(3) xor hash_input(7) xor hash_input(10) xor hash_input(11) xor hash_input(13) xor hash_input(14) xor hash_input(16) xor hash_input(18) xor hash_input(20) xor hash_input(31) xor hash_input(33) xor hash_input(34) xor hash_input(38) xor hash_input(41) xor hash_input(42) xor hash_input(44) xor hash_input(45) xor hash_input(47) xor hash_input(49) xor hash_input(51) xor hash_input(62) xor hash_input(64) xor hash_input(65) xor hash_input(69) xor hash_input(72) xor hash_input(73) xor hash_input(75) xor hash_input(76) xor hash_input(78) xor hash_input(80) xor hash_input(82) xor hash_input(93) xor hash_input(95) xor hash_input(96) xor hash_input(100) xor hash_input(103) ; 
	hash_output(1) <= hash_input(1) xor hash_input(3) xor hash_input(4) xor hash_input(8) xor hash_input(11) xor hash_input(12) xor hash_input(14) xor hash_input(15) xor hash_input(17) xor hash_input(19) xor hash_input(21) xor hash_input(32) xor hash_input(34) xor hash_input(35) xor hash_input(39) xor hash_input(42) xor hash_input(43) xor hash_input(45) xor hash_input(46) xor hash_input(48) xor hash_input(50) xor hash_input(52) xor hash_input(63) xor hash_input(65) xor hash_input(66) xor hash_input(70) xor hash_input(73) xor hash_input(74) xor hash_input(76) xor hash_input(77) xor hash_input(79) xor hash_input(81) xor hash_input(83) xor hash_input(94) xor hash_input(96) xor hash_input(97) xor hash_input(101) ; 
	hash_output(2) <= hash_input(0) xor hash_input(3) xor hash_input(4) xor hash_input(5) xor hash_input(7) xor hash_input(9) xor hash_input(10) xor hash_input(11) xor hash_input(12) xor hash_input(14) xor hash_input(15) xor hash_input(22) xor hash_input(31) xor hash_input(34) xor hash_input(35) xor hash_input(36) xor hash_input(38) xor hash_input(40) xor hash_input(41) xor hash_input(42) xor hash_input(43) xor hash_input(45) xor hash_input(46) xor hash_input(53) xor hash_input(62) xor hash_input(65) xor hash_input(66) xor hash_input(67) xor hash_input(69) xor hash_input(71) xor hash_input(72) xor hash_input(73) xor hash_input(74) xor hash_input(76) xor hash_input(77) xor hash_input(84) xor hash_input(93) xor hash_input(96) xor hash_input(97) xor hash_input(98) xor hash_input(100) xor hash_input(102) xor hash_input(103) ; 
	hash_output(3) <= hash_input(1) xor hash_input(4) xor hash_input(5) xor hash_input(6) xor hash_input(8) xor hash_input(10) xor hash_input(11) xor hash_input(12) xor hash_input(13) xor hash_input(15) xor hash_input(16) xor hash_input(23) xor hash_input(32) xor hash_input(35) xor hash_input(36) xor hash_input(37) xor hash_input(39) xor hash_input(41) xor hash_input(42) xor hash_input(43) xor hash_input(44) xor hash_input(46) xor hash_input(47) xor hash_input(54) xor hash_input(63) xor hash_input(66) xor hash_input(67) xor hash_input(68) xor hash_input(70) xor hash_input(72) xor hash_input(73) xor hash_input(74) xor hash_input(75) xor hash_input(77) xor hash_input(78) xor hash_input(85) xor hash_input(94) xor hash_input(97) xor hash_input(98) xor hash_input(99) xor hash_input(101) xor hash_input(103) ; 
	hash_output(4) <= hash_input(2) xor hash_input(5) xor hash_input(6) xor hash_input(7) xor hash_input(9) xor hash_input(11) xor hash_input(12) xor hash_input(13) xor hash_input(14) xor hash_input(16) xor hash_input(17) xor hash_input(24) xor hash_input(33) xor hash_input(36) xor hash_input(37) xor hash_input(38) xor hash_input(40) xor hash_input(42) xor hash_input(43) xor hash_input(44) xor hash_input(45) xor hash_input(47) xor hash_input(48) xor hash_input(55) xor hash_input(64) xor hash_input(67) xor hash_input(68) xor hash_input(69) xor hash_input(71) xor hash_input(73) xor hash_input(74) xor hash_input(75) xor hash_input(76) xor hash_input(78) xor hash_input(79) xor hash_input(86) xor hash_input(95) xor hash_input(98) xor hash_input(99) xor hash_input(100) xor hash_input(102) ; 
	hash_output(5) <= hash_input(3) xor hash_input(6) xor hash_input(7) xor hash_input(8) xor hash_input(10) xor hash_input(12) xor hash_input(13) xor hash_input(14) xor hash_input(15) xor hash_input(17) xor hash_input(18) xor hash_input(25) xor hash_input(34) xor hash_input(37) xor hash_input(38) xor hash_input(39) xor hash_input(41) xor hash_input(43) xor hash_input(44) xor hash_input(45) xor hash_input(46) xor hash_input(48) xor hash_input(49) xor hash_input(56) xor hash_input(65) xor hash_input(68) xor hash_input(69) xor hash_input(70) xor hash_input(72) xor hash_input(74) xor hash_input(75) xor hash_input(76) xor hash_input(77) xor hash_input(79) xor hash_input(80) xor hash_input(87) xor hash_input(96) xor hash_input(99) xor hash_input(100) xor hash_input(101) xor hash_input(103) ; 
	hash_output(6) <= hash_input(4) xor hash_input(7) xor hash_input(8) xor hash_input(9) xor hash_input(11) xor hash_input(13) xor hash_input(14) xor hash_input(15) xor hash_input(16) xor hash_input(18) xor hash_input(19) xor hash_input(26) xor hash_input(35) xor hash_input(38) xor hash_input(39) xor hash_input(40) xor hash_input(42) xor hash_input(44) xor hash_input(45) xor hash_input(46) xor hash_input(47) xor hash_input(49) xor hash_input(50) xor hash_input(57) xor hash_input(66) xor hash_input(69) xor hash_input(70) xor hash_input(71) xor hash_input(73) xor hash_input(75) xor hash_input(76) xor hash_input(77) xor hash_input(78) xor hash_input(80) xor hash_input(81) xor hash_input(88) xor hash_input(97) xor hash_input(100) xor hash_input(101) xor hash_input(102) ; 
	hash_output(7) <= hash_input(0) xor hash_input(2) xor hash_input(3) xor hash_input(5) xor hash_input(7) xor hash_input(8) xor hash_input(9) xor hash_input(11) xor hash_input(12) xor hash_input(13) xor hash_input(15) xor hash_input(17) xor hash_input(18) xor hash_input(19) xor hash_input(27) xor hash_input(31) xor hash_input(33) xor hash_input(34) xor hash_input(36) xor hash_input(38) xor hash_input(39) xor hash_input(40) xor hash_input(42) xor hash_input(43) xor hash_input(44) xor hash_input(46) xor hash_input(48) xor hash_input(49) xor hash_input(50) xor hash_input(58) xor hash_input(62) xor hash_input(64) xor hash_input(65) xor hash_input(67) xor hash_input(69) xor hash_input(70) xor hash_input(71) xor hash_input(73) xor hash_input(74) xor hash_input(75) xor hash_input(77) xor hash_input(79) xor hash_input(80) xor hash_input(81) xor hash_input(89) xor hash_input(93) xor hash_input(95) xor hash_input(96) xor hash_input(98) xor hash_input(100) xor hash_input(101) xor hash_input(102) ; 
	hash_output(8) <= hash_input(0) xor hash_input(1) xor hash_input(2) xor hash_input(4) xor hash_input(6) xor hash_input(7) xor hash_input(8) xor hash_input(9) xor hash_input(11) xor hash_input(12) xor hash_input(19) xor hash_input(28) xor hash_input(31) xor hash_input(32) xor hash_input(33) xor hash_input(35) xor hash_input(37) xor hash_input(38) xor hash_input(39) xor hash_input(40) xor hash_input(42) xor hash_input(43) xor hash_input(50) xor hash_input(59) xor hash_input(62) xor hash_input(63) xor hash_input(64) xor hash_input(66) xor hash_input(68) xor hash_input(69) xor hash_input(70) xor hash_input(71) xor hash_input(73) xor hash_input(74) xor hash_input(81) xor hash_input(90) xor hash_input(93) xor hash_input(94) xor hash_input(95) xor hash_input(97) xor hash_input(99) xor hash_input(100) xor hash_input(101) xor hash_input(102) ; 
	hash_output(9) <= hash_input(0) xor hash_input(1) xor hash_input(5) xor hash_input(8) xor hash_input(9) xor hash_input(11) xor hash_input(12) xor hash_input(14) xor hash_input(16) xor hash_input(18) xor hash_input(29) xor hash_input(31) xor hash_input(32) xor hash_input(36) xor hash_input(39) xor hash_input(40) xor hash_input(42) xor hash_input(43) xor hash_input(45) xor hash_input(47) xor hash_input(49) xor hash_input(60) xor hash_input(62) xor hash_input(63) xor hash_input(67) xor hash_input(70) xor hash_input(71) xor hash_input(73) xor hash_input(74) xor hash_input(76) xor hash_input(78) xor hash_input(80) xor hash_input(91) xor hash_input(93) xor hash_input(94) xor hash_input(98) xor hash_input(101) xor hash_input(102) ; 
	hash_output(10) <= hash_input(1) xor hash_input(2) xor hash_input(6) xor hash_input(9) xor hash_input(10) xor hash_input(12) xor hash_input(13) xor hash_input(15) xor hash_input(17) xor hash_input(19) xor hash_input(30) xor hash_input(32) xor hash_input(33) xor hash_input(37) xor hash_input(40) xor hash_input(41) xor hash_input(43) xor hash_input(44) xor hash_input(46) xor hash_input(48) xor hash_input(50) xor hash_input(61) xor hash_input(63) xor hash_input(64) xor hash_input(68) xor hash_input(71) xor hash_input(72) xor hash_input(74) xor hash_input(75) xor hash_input(77) xor hash_input(79) xor hash_input(81) xor hash_input(92) xor hash_input(94) xor hash_input(95) xor hash_input(99) xor hash_input(102) xor hash_input(103) ; 
end generate;
	
hash_funct_10bits: if(OUTPUT_WIDTH = 10) generate
	hash_output(0) <= hash_input(0) xor hash_input(1) xor hash_input(2) xor hash_input(3) xor hash_input(4) xor hash_input(9) xor hash_input(15) xor hash_input(16) xor hash_input(17) xor hash_input(19) xor hash_input(23) xor hash_input(24) xor hash_input(27) xor hash_input(28) xor hash_input(30) xor hash_input(31) xor hash_input(32) xor hash_input(33) xor hash_input(34) xor hash_input(36) xor hash_input(37) xor hash_input(39) xor hash_input(41) xor hash_input(42) xor hash_input(46) xor hash_input(49) xor hash_input(51) xor hash_input(52) xor hash_input(53) xor hash_input(58) xor hash_input(59) xor hash_input(65) xor hash_input(66) xor hash_input(69) xor hash_input(72) xor hash_input(73) xor hash_input(74) xor hash_input(76) xor hash_input(78) xor hash_input(80) xor hash_input(81) xor hash_input(83) xor hash_input(84) xor hash_input(85) xor hash_input(89) xor hash_input(90) xor hash_input(91) xor hash_input(94) xor hash_input(97) xor hash_input(99) xor hash_input(101) ; 
	hash_output(1) <= hash_input(0) xor hash_input(5) xor hash_input(9) xor hash_input(10) xor hash_input(15) xor hash_input(18) xor hash_input(19) xor hash_input(20) xor hash_input(23) xor hash_input(25) xor hash_input(27) xor hash_input(29) xor hash_input(30) xor hash_input(35) xor hash_input(36) xor hash_input(38) xor hash_input(39) xor hash_input(40) xor hash_input(41) xor hash_input(43) xor hash_input(46) xor hash_input(47) xor hash_input(49) xor hash_input(50) xor hash_input(51) xor hash_input(54) xor hash_input(58) xor hash_input(60) xor hash_input(65) xor hash_input(67) xor hash_input(69) xor hash_input(70) xor hash_input(72) xor hash_input(75) xor hash_input(76) xor hash_input(77) xor hash_input(78) xor hash_input(79) xor hash_input(80) xor hash_input(82) xor hash_input(83) xor hash_input(86) xor hash_input(89) xor hash_input(92) xor hash_input(94) xor hash_input(95) xor hash_input(97) xor hash_input(98) xor hash_input(99) xor hash_input(100) xor hash_input(101) xor hash_input(102) ; 
	hash_output(2) <= hash_input(1) xor hash_input(6) xor hash_input(10) xor hash_input(11) xor hash_input(16) xor hash_input(19) xor hash_input(20) xor hash_input(21) xor hash_input(24) xor hash_input(26) xor hash_input(28) xor hash_input(30) xor hash_input(31) xor hash_input(36) xor hash_input(37) xor hash_input(39) xor hash_input(40) xor hash_input(41) xor hash_input(42) xor hash_input(44) xor hash_input(47) xor hash_input(48) xor hash_input(50) xor hash_input(51) xor hash_input(52) xor hash_input(55) xor hash_input(59) xor hash_input(61) xor hash_input(66) xor hash_input(68) xor hash_input(70) xor hash_input(71) xor hash_input(73) xor hash_input(76) xor hash_input(77) xor hash_input(78) xor hash_input(79) xor hash_input(80) xor hash_input(81) xor hash_input(83) xor hash_input(84) xor hash_input(87) xor hash_input(90) xor hash_input(93) xor hash_input(95) xor hash_input(96) xor hash_input(98) xor hash_input(99) xor hash_input(100) xor hash_input(101) xor hash_input(102) xor hash_input(103) ; 
	hash_output(3) <= hash_input(2) xor hash_input(7) xor hash_input(11) xor hash_input(12) xor hash_input(17) xor hash_input(20) xor hash_input(21) xor hash_input(22) xor hash_input(25) xor hash_input(27) xor hash_input(29) xor hash_input(31) xor hash_input(32) xor hash_input(37) xor hash_input(38) xor hash_input(40) xor hash_input(41) xor hash_input(42) xor hash_input(43) xor hash_input(45) xor hash_input(48) xor hash_input(49) xor hash_input(51) xor hash_input(52) xor hash_input(53) xor hash_input(56) xor hash_input(60) xor hash_input(62) xor hash_input(67) xor hash_input(69) xor hash_input(71) xor hash_input(72) xor hash_input(74) xor hash_input(77) xor hash_input(78) xor hash_input(79) xor hash_input(80) xor hash_input(81) xor hash_input(82) xor hash_input(84) xor hash_input(85) xor hash_input(88) xor hash_input(91) xor hash_input(94) xor hash_input(96) xor hash_input(97) xor hash_input(99) xor hash_input(100) xor hash_input(101) xor hash_input(102) xor hash_input(103) ; 
	hash_output(4) <= hash_input(0) xor hash_input(1) xor hash_input(2) xor hash_input(4) xor hash_input(8) xor hash_input(9) xor hash_input(12) xor hash_input(13) xor hash_input(15) xor hash_input(16) xor hash_input(17) xor hash_input(18) xor hash_input(19) xor hash_input(21) xor hash_input(22) xor hash_input(24) xor hash_input(26) xor hash_input(27) xor hash_input(31) xor hash_input(34) xor hash_input(36) xor hash_input(37) xor hash_input(38) xor hash_input(43) xor hash_input(44) xor hash_input(50) xor hash_input(51) xor hash_input(54) xor hash_input(57) xor hash_input(58) xor hash_input(59) xor hash_input(61) xor hash_input(63) xor hash_input(65) xor hash_input(66) xor hash_input(68) xor hash_input(69) xor hash_input(70) xor hash_input(74) xor hash_input(75) xor hash_input(76) xor hash_input(79) xor hash_input(82) xor hash_input(84) xor hash_input(86) xor hash_input(90) xor hash_input(91) xor hash_input(92) xor hash_input(94) xor hash_input(95) xor hash_input(98) xor hash_input(99) xor hash_input(100) xor hash_input(102) xor hash_input(103) ; 
	hash_output(5) <= hash_input(0) xor hash_input(4) xor hash_input(5) xor hash_input(10) xor hash_input(13) xor hash_input(14) xor hash_input(15) xor hash_input(18) xor hash_input(20) xor hash_input(22) xor hash_input(24) xor hash_input(25) xor hash_input(30) xor hash_input(31) xor hash_input(33) xor hash_input(34) xor hash_input(35) xor hash_input(36) xor hash_input(38) xor hash_input(41) xor hash_input(42) xor hash_input(44) xor hash_input(45) xor hash_input(46) xor hash_input(49) xor hash_input(53) xor hash_input(55) xor hash_input(60) xor hash_input(62) xor hash_input(64) xor hash_input(65) xor hash_input(67) xor hash_input(70) xor hash_input(71) xor hash_input(72) xor hash_input(73) xor hash_input(74) xor hash_input(75) xor hash_input(77) xor hash_input(78) xor hash_input(81) xor hash_input(84) xor hash_input(87) xor hash_input(89) xor hash_input(90) xor hash_input(92) xor hash_input(93) xor hash_input(94) xor hash_input(95) xor hash_input(96) xor hash_input(97) xor hash_input(100) xor hash_input(103) ; 
	hash_output(6) <= hash_input(1) xor hash_input(5) xor hash_input(6) xor hash_input(11) xor hash_input(14) xor hash_input(15) xor hash_input(16) xor hash_input(19) xor hash_input(21) xor hash_input(23) xor hash_input(25) xor hash_input(26) xor hash_input(31) xor hash_input(32) xor hash_input(34) xor hash_input(35) xor hash_input(36) xor hash_input(37) xor hash_input(39) xor hash_input(42) xor hash_input(43) xor hash_input(45) xor hash_input(46) xor hash_input(47) xor hash_input(50) xor hash_input(54) xor hash_input(56) xor hash_input(61) xor hash_input(63) xor hash_input(65) xor hash_input(66) xor hash_input(68) xor hash_input(71) xor hash_input(72) xor hash_input(73) xor hash_input(74) xor hash_input(75) xor hash_input(76) xor hash_input(78) xor hash_input(79) xor hash_input(82) xor hash_input(85) xor hash_input(88) xor hash_input(90) xor hash_input(91) xor hash_input(93) xor hash_input(94) xor hash_input(95) xor hash_input(96) xor hash_input(97) xor hash_input(98) xor hash_input(101) ; 
	hash_output(7) <= hash_input(2) xor hash_input(6) xor hash_input(7) xor hash_input(12) xor hash_input(15) xor hash_input(16) xor hash_input(17) xor hash_input(20) xor hash_input(22) xor hash_input(24) xor hash_input(26) xor hash_input(27) xor hash_input(32) xor hash_input(33) xor hash_input(35) xor hash_input(36) xor hash_input(37) xor hash_input(38) xor hash_input(40) xor hash_input(43) xor hash_input(44) xor hash_input(46) xor hash_input(47) xor hash_input(48) xor hash_input(51) xor hash_input(55) xor hash_input(57) xor hash_input(62) xor hash_input(64) xor hash_input(66) xor hash_input(67) xor hash_input(69) xor hash_input(72) xor hash_input(73) xor hash_input(74) xor hash_input(75) xor hash_input(76) xor hash_input(77) xor hash_input(79) xor hash_input(80) xor hash_input(83) xor hash_input(86) xor hash_input(89) xor hash_input(91) xor hash_input(92) xor hash_input(94) xor hash_input(95) xor hash_input(96) xor hash_input(97) xor hash_input(98) xor hash_input(99) xor hash_input(102) ; 
	hash_output(8) <= hash_input(3) xor hash_input(7) xor hash_input(8) xor hash_input(13) xor hash_input(16) xor hash_input(17) xor hash_input(18) xor hash_input(21) xor hash_input(23) xor hash_input(25) xor hash_input(27) xor hash_input(28) xor hash_input(33) xor hash_input(34) xor hash_input(36) xor hash_input(37) xor hash_input(38) xor hash_input(39) xor hash_input(41) xor hash_input(44) xor hash_input(45) xor hash_input(47) xor hash_input(48) xor hash_input(49) xor hash_input(52) xor hash_input(56) xor hash_input(58) xor hash_input(63) xor hash_input(65) xor hash_input(67) xor hash_input(68) xor hash_input(70) xor hash_input(73) xor hash_input(74) xor hash_input(75) xor hash_input(76) xor hash_input(77) xor hash_input(78) xor hash_input(80) xor hash_input(81) xor hash_input(84) xor hash_input(87) xor hash_input(90) xor hash_input(92) xor hash_input(93) xor hash_input(95) xor hash_input(96) xor hash_input(97) xor hash_input(98) xor hash_input(99) xor hash_input(100) xor hash_input(103) ; 
	hash_output(9) <= hash_input(0) xor hash_input(1) xor hash_input(2) xor hash_input(3) xor hash_input(8) xor hash_input(14) xor hash_input(15) xor hash_input(16) xor hash_input(18) xor hash_input(22) xor hash_input(23) xor hash_input(26) xor hash_input(27) xor hash_input(29) xor hash_input(30) xor hash_input(31) xor hash_input(32) xor hash_input(33) xor hash_input(35) xor hash_input(36) xor hash_input(38) xor hash_input(40) xor hash_input(41) xor hash_input(45) xor hash_input(48) xor hash_input(50) xor hash_input(51) xor hash_input(52) xor hash_input(57) xor hash_input(58) xor hash_input(64) xor hash_input(65) xor hash_input(68) xor hash_input(71) xor hash_input(72) xor hash_input(73) xor hash_input(75) xor hash_input(77) xor hash_input(79) xor hash_input(80) xor hash_input(82) xor hash_input(83) xor hash_input(84) xor hash_input(88) xor hash_input(89) xor hash_input(90) xor hash_input(93) xor hash_input(96) xor hash_input(98) xor hash_input(100) ; 	
end generate;

end architecture hash_function_arch;

