XlxV64EB    5185    1230I��P=`�O緼����ʙ�T����7ڻ��^�p�*���h1-�rc�s�
���%w[�>m�;�.��Bl��%�ii�q��nKo��@gJ_�ƪK��w
��A��%8���n�^5��QT�˪}^b!�Mʅ��3��/��S ��Vw�Ǫ �w��	��4p�a�O���R* �;�0}*��ۤ���>��d'��/-+z�E�;�3�Y���}�a��V�F�T��vHD��=��H_&��_<������4�i7��M��f�-KP��P8�^��u
�{����Nc}�:Bڵ�XJA��ڬ-�FޅX�/J�𓘕o�Y	�s��.$�M+�|$LƆQ��R���ᘅ��~���8vR����xr���+1��%�k�{?f�@�bY�����Α�����R��1z��fU=��1���$Ę?f�QMdt��g���S&��4�U*�h26��s]�Mx�����J������� 6�]�&�5�֤<ׁ�@�]�ʩ}	җK�~=,�n+3]� ��[/��yl���f`gz���� �B�Q8U�^f��0d��<��?ft(h�i# z��a�V�P*H:(ܣ�*7`�VQ�Q�\�o��NLzA���J3o��	t"��g�^��j���2�{W�UΏ��˕ e;sK>/u�9L6 �Avgъ�f�p~�F��@|�������[t*�6�x�1�Q��i2����sM57w�:6���n&�*�f�B06_���C�>��c�r��^�*�� _0�L_��B��ѐ�/ .�k��پ�T��%:0H�8[јh[�2g�=����8T(�Ժ��C�I�R5v|�|v��&�z�eF��5ݡ���:;�X���G�cU��^�[�&D^��VK�cB�~CN5�h���QSa{����_�iE90�r�W��J`]�`d?�Ku$<�N<���u5k<�_(^�����FER���N�o(E�߈=��tQ�وI{ &Ή� ���(��rî�&l9^��8ֻ�h72��N@���ͯw��!��䘧��]�I��]?L�[���	h��tC}�w4��v�f_4B⿡�	ش	��U��%yYͥ�b��ֹ�YH�����2%�L��Cv��孬BԞ�u<'����]�v,�i<���.�Y�!s�Z�5�%�����H��W��0�J͟AJE:P�2�՟cd�m���C��Ţ=!0�Y�ua-؀�y�m���=�MP�
dđ��qR(����_�_>}�O��S��K�gs�Hх<�J�ʌ��y�r���sr�V��G�>��;#Q���Z\YWN�P!E'޷��L�����2���i�id�-�b�|!���$uz��`��S?g	�·��Ra��� ����1�*�G	�g��$c���%DGYu�q��\���R#�-z�c�jcQ\}(yC5�f�Dc���R���?�aL]��Su�y��(�Z�7Z��E(=�_�ܙx�^V�d�����{�"t%�g�n�?���
�=1⌣��Z��/5����=ߋ>:Y�N�f��'75K緍B���ǐ
���w����N��Q�H���[�Z�<~�N)Q�ڢ�9���SİD��K�&eǸ*o����/+	-�pTh��IR-*6,BTzB��{[��/R��c� YC����[0�,���PזB>�[����O��Z��,���~N��Q���Gc�_��� e�`x�[L�n�E�XE�&��$y��
�?�fG�Ϥp�\-�����f+�̄�e u&:�'�5p�*�A�o��D^p�,焒�ȚP��P3q�uC��7�T�t���a�:N�K���X��UBmw���8I<Q�:��F��5���m����U~d�@��l˖�
��~��	iEk��|p[r'ɏ"Eڣ�Vn0b� ~7'f�R���M����lie��l����(�ư*�lZ��[��/�T�@��Rē�k8�3���Z�S�GУ�6�끢��n�R��;�g�ܓ
�'m��\C�ޛ������F�-�����e�7�2��t�G
�.��O�������c��V�����w�4�,��+�a�k�6p�T��t����dzB�Aᅧ0tH6w�&��e�^72�,�Τ5YF��ux�+���A��.���'2PI{��O�����6�s�0AbB}�� 	G%��ą+D������h�G����[�"#���C��p�7E�|�����j��]+o)*���J�!40u�}�]v��ZOY�/�jmk_6N�� �~�����õG:@��nڊKN�7���eC�v+��˯����$r4�sK]�j�i�m(�/}���[�+�$���j�yK�7�]z��QS�tL�,�Qe-�r�~t=C��&�U�}��yB�5$+��	|�3���d���(馄m1K���>��z���ԿN�����N �N�Ѿu���t�v����F���f�b�I�K[N2 ����mr�l���`-���+�7��k�F�c�"fF;��Z�C��O]y�1��V9��%Ζ $Q� 5jR�hʥ1\��HL?pK�@� ��� �;��pŻk���
�6W��EV�~B?��h[����+�/��~��E���O�����kI���N�6�p5�NkK��:H���S��Nx��,��[�{�JK�:g&���:�-2���v#(��Z�k�Rf֤�����BF	�:ʓ���	��1��5@�(��w�M�#D�:�9�NeL��!I˚�lD�.����d���E-H���Cdb�1����֣���)p�b5ފu���ό�٤φB�ڜ�3���|b���y���e+6넂��%p������ư�ߌP>T��Q`ؐ�J�ƙdn�މ�D�,]C�pZ��(���#��`�A;uh;=t?Aۚ���B���G�[r?��j��8�Q�B���5��z����&V��k�3�Y��P,����}r8����5 �<�o[������c�Ƃ����FȒ0Â��2�����z�ݺk�C���:]Bͤ�����ʗq'Aڼh���X����_��
����M훾��t��{ =0��4�}S������Ļ`�"�|"�ZaɃl ���HX��I�3*a�{F�F�T�C`4��G=DA/��NE#�����	����M�Z�DU�y��ft����1�2�hB����_:Ͼ�T[���C����.U/�/lR���'��ޏ@�e�w������2W>�|�p���z��1-$�x~
Q���T�Ƈ��I�@��FX�UV�ޯ�Rjv?��	�/�h���J�j�z_���'���Z�$���Wu��9Wˇ����	�E<�̛!�1%tH��g%�¾|CF_q��#$m7#m��< �7�#e���@�V� �nH�r�z�+�g�ʋ1�(�\��_���հ~ԭ1H���?���-�`�_?Z6��Jğ)�$���,�- �+	ˍ��=gȝ�4��~�6��P��H�ZA�N=B�<
k�E����fA#G���h�ѺY�q�E8%������T=`��·)����	ߜ!H�&�O��؇�4_�9	֍�=�;��н���d�wXPD�xj-��W6J���v��,ܿ	NŘ,��~z� S�l���	.�xHuG챐wg��?N��Ȕ6̵@��Uh��o�7u1�3�$�mX;y<;�$!D ♶�,l��p��[��Χ�|�1#>.3?B4����T޳=�$��sS|�Q5+�����#�f��˃i#S|t�H�W���)���'�3������CX� ��A&4��GOT]�K�ٛ���arS����,yJML���#[��)ۤC`�c�[�5,	y!\o�M�⇃sK�\�߹���ח[B�~8"T٪�rș\�^3`klC;�'ަ��x%nl!u^��5�
�����Tg�P ;@��������Z���4�[
EN�oKp�eaG�`5�:�v��!� BQ��t���LLH[s�����{�1��Q��tٕ=#������y�q$���} ��1fTse�D�Q��������\�-Q~��3Ԡ.�yjG�3�����J�3T1W#	��4��\E5]�q�CFײ��K��y�̬s�Mz�v����?�n�:���x�LȧqnE����p�K��N�}d�a�V��u���
�C��v�0|Ok�i��(����I>r� ;�*��Ӽ����ܭq>�c;�1�>��Jb>�\��H��pS1גN�vei���������`��q�p�[,'/���i�E�=�I��Z�Y�SC��#��PAnr6�P�]�S��̿�7��P<`��c�7N,+l3C꥾��kלENk��lm��ь�s�Ѣ��j�L�_��B��]Z���1�y�oQ-JQ�:�.o����7����̠�SD�>�`����w�B9ѩX�p���n�c�Z,r�R+�R��El8�&�V�N��M����6H����H/i��y)b���u�ܥ`k�R)j:`�W̅�s��<�ؤ��+��{cA��q˺ɜ��.	b�t�#�}e�S��|܃2�tV}��E4�]^l�#����Jl��(�n���-h��!:ဗ�