XlxV64EB    17fc     9b0��b�O�� ��z���;#_1DC�B�����hN��W��R��\o�C�0%���C�E�2��_1d=�y�����RD�GKB��ż$I�J�R�^Fyp���x���R�2�;!�d�$��"��a�09��P�
P�Eq��6,j@��mI��;k+�~����V�KG���X��P��*{�Y��c���P)A�'�Tg�ic���4+�[�$65T�y�n�,�5E`�w��ȉ>='�F�uuoh�������������oZ���M�g�ώج�7'Ac'G��!�e�A�X$���0
\��J�u}�phWG�Yg�4Ͼ!I��]��׋���1ʻR;�_ThPr�4O��3UP��pb���36ק��/���p�tR(�z�Hs�2b�F�y3<�O��x�v�QFA��u�%����K�f�X<����Fd����5�8�En$�Y����ÏY]�@bumۼ����&�ghl־��Ge���������ؗ	����v[%6��8�@���7�1n�
�� �ڔ�9X�:��┩�f��B�i���9	J��l*�"@g]�����6�@�I	���J)EO�':T���]`rSNO�w4�kڮ��aն�����FC8&e?N�/�2�kDX�?�V�{�y���n�%��3L{�[�O�E!>��L���G,� �J��͆��d�B=�}�{�1C����bD����&W}�(�e~m�X��H�]�F�Ǹ7��<p%�v�&tuiA� ��7+�D�ba�8j��9�����sZ�b|����L5F>���=��l$6l��dѪ��8��QC_�$�#��,lѵ�i.t=������������i����ɾc��9�9Hz�l$q��?�L�/��,���A2¾�������V57����^�>!�OK ���7�b��0���gD̞��2�s�D��2Z-�V�輌f�P�����A�~#{@���J)�~��(�����+��,ʇ��T a����w��,�U����K"*2��;��^)��)Y {d�ƹ�GV:^�v?�?���˷�!�D9˵8�E���9_1��Aam1M��=:�zo}�Z�7�1S^��vbK6B&� GZ[��"&�;�խٜ�d�30���K��3�����j��\��s�E�[�Q�m���!�~������'넙��<w�&?GKp7������ s
5���O]��� �M�S�CϤ�{3	�C;Y�ʲ�t ��*��.F�i�Qz yw^n1t�+<�4��M;?
�a��@��3.Y 5�CbK_�Tj��A0�r�WN[�׾_��|�	'�+�N��fg�������8	ۈjn�v���C�ǀ�%�P`�ՃT�#��z��m �T�(�n�Y�Ɲe��٨A
m͉�fm^�r=��ϾF=�+���L� � �kI$
���{�tH؀
���'�U�>:�Jgl�cm~��w����ְ�.9�؞���1��LS�0F��x׶p�-:�Ê��P$�C9(y ݳw�y`���8���	|�C�@�6��%8���ü�Rg�=d��D!G9-Ra�0N实ᨗ���ǝ��U[���<�IC���^s��WvqA�M�H�m"8P�S�ڒN.��`gHm5
�j
���kq�A���rFؼ3�CRB �i�s��;�ӂy��io�}�^ߔ�Iy����ϐX2���8���|d2s�<~�կ��o�=
h	�Z�R�.� t��W�x�+Vo�\�N��֐џ��U8�1Z�"˅l.!nqCn:����	nƽ�0@u�}%��I�!����>1����V	��"�U�=JؙG��7���B/�5ļ_�5�gD�>�3�A��M�"���<q�SC��j-�?:���������ʆ�s��ˉ%�k����Y�S�}�>$$eA8}RߌV��/D	���VY�d��/	��9?D�:=?eN=�#\�u]tl Ta���=C�"�Ńc�Wˮ�)��:����R��Bʶh��+����f�ʺ��+|�'?��yūhn��벟M�)L+/�n��@���0�����#� &1C]�2qCPNn�P�Q��	��Ӓ�y�#c�3
R����s���b��	�9�ߗ�t`@ߍ�e9��Y�QU�dSZ��x�4��\5�R�4�i;��l"��C3�7my�u�0�K�`�OE��
A�F����?��L[���g4"�>�Q5p#�"b��ie��%�|\k�J��e�_<��F� ���]*Vx#��Y[J+�w�_^gkKQ�l8���D�l{q��Y5���z��Ndsn_Z�F�
��Q\�+�r
�<y&A�|C�b�ֻϷ�O	ht�3�m����R4���H*f0���:7ETq����$[%:�LQ��Ks_��O�X+��[�����u�ŴG��H��?H~��gl�:j�?<{��wt�r�l�1=�<�H&��9�K�'\�.��N:	T֔g��y|�0L�Mo�̲�