XlxV64EB    2599     b40�.U)Qp�iD4pVCu��"n� ��O��H�:L���ǘ����S=��1���
3qfO�`��ҥL̀��l�ʅ���ԝ7��|����"m�2�y1iP�;i�w��1�Y��N�02�!#_l,p���Qs$ҎyÊB�hi|��
+Dw�4��8�����`�Z1:���:ؔ�L���Yj��5f��i���s�΢]W���q���=IA�ƶڠ�庄�|؀�!V�3�m���s�c����
�+OlEyӝ����8�T�ƥhߐ���1g�.�#�����X�:==o�P�Pw�E	�z0G*���`/ɬ>Еx��
��n��~;�Ӛ��䄅�G���{��{�׌�8��T�݋�Ā�cB�3r�6��^X�N?٢�-��l�!��47%O���_�.܉,�� ��>`~h��C�a��;]̝=']��J7�j�v,�.v�;+8]
т�����6�Ҕ�b.F�e���W�ϓt(��_v��^_����6� �d:��Cr�=l/T'�j��㕾���ng�xGi���^��� G�1��o5�s�(;W�,V�����i���)τ$O�jL�-�&%�,�Lz߫~��ɭ���D@Q�0��m�z,��<�謐<�zч�.%%(���+�:v/�](g��_���̗��H�ri���������ek�`�؁�N
��^,:���PT�9����DG��l4��zKX�Y� ���qK�����B}�� S?����[�%6�̅벣 1b�R�H_7��Ǝ�`��z�l���uL3|���Oݱ�R�R�)��"��}����Ӿ1w1.h��س�'霯ז�Nb R�,�Qr ix�� ����u!�eU��UC����7O������&�@z��[�e3DV�r�B����x��j�f͡wq�k�I�� �I�5�L��f�������s���t!q�T���Y�h��C�g�S-��+r>P.,��T�&���Z0���������0P��<�-y��}!�Mf�>Q��0W.�i�K��h�7f��� u�J��a��nj9�U�8�#�Lo�&eϵ�R~/�1�+�VBֵ���n�b�L���
-f[/9���f�n�\��wN���S��[֋c^	:�L�h5}��+8������f����]��wIQ'G�*M�D*9�"�b�bSƺw@s�M��P�^����	�X��3�����<rnM�������Gרt{
�t�`&���du�/�?o���@��1�B��ln�=���smn�;�Ğ ���ibw��px�1�*!-��=��Q�jO�|��;])$����zf�D��3���Wƿ#ax�R�0�1a)���Q=8�,)��(�?�G��-ˀN�������ʦ��_��O^������јCk�o#b��U��S���Rn)��g�W���m<��E[��a4Pn7ߝ	�\t5��㿮I�@��	���B���4�I�����֩w�Z��
���Q(#c0���se���]i�K.�9Ola�)f��d�ސ��@t���kE(��NɽlO�y %�-�y�'��Ϻ��z�2i��@��M�,��=�d��&��1�:���_�S7~�y�W9bK��uIH�᭨���f��}��:x$Z����l~�.���}���.s�S+�'��t�:�^�4Y��d�f�e/.v�0c|Ι�d�'�}\Y�"��Q�>r4U��9L�� /�}4��J�����BԶ=�L�4g�r\���	�$텱*���Ћ9]�z�,��L����*�X�����Sp�Ć;�8�$����fuVH3L�D�ZP0��B)���,�Ll/�F՝�Z���� #+�lE������z�,�Gl�*����� f~4FWA(rrW��l&wI�f���'c+5�K�v=�0�R)V=����DML���#�=�E�nw/�K����iս�����q�#��4�}����V�@���ɟ��X����xzDU>jѸC�� ��]��r�~r�i�S��s�<z7$�68f�b�^��f�GSm���=�� �_���V�Ye�=fɀN��/٭QU����%<Y�C�m�Zr�p���.w�>Q�Xc#7����R��IMDiʹ1�ߞ�:�\��:�H�R+/�}"�5�W��8��XࡋLo`�I�k)����&���ӯ�O[:R��1)����-,�f�G��&j�Q��Ih8p��w�L>w�Gl����B�E��'���*�Q_�Gq�q�$*��t+��8��)�>��[L������R�*�`815<�<*���k	x)'��%o$X����D
�F:�9ϐ*u��+'�����1�ן���!��[e&R�Y=��� u�P�?^/�������J_���4A�vQˀ���i���?L��>�i�QӋ�KD��� 3����c>3�ޭnN�� ���,��$�����bӌ�w��A��x��.�%�M�7d�=�m|S ��ީv�ySe1!�9���Dtc&����+�	SN��z��ǔ�܂=�Z׺@򰐡sFZ��=��<2\�"�7>F\Vodo_,�Q���&�9uc�赿�i�?V;��N����_xeAN�\1;�$��]~P��Ӑ���NU�_7Y�ȭ]���[[CU@��y�����^��6��ǒ�қ���2�Θ�������́@G�h>2�X2	{���j��戌�&_�����k�o�;�� j�Em\��t�=(o���P6P������^�0F�ca���:�:Y�˵.�gh��>����B��˖��{7=Ki�{�m�������y��IS<4�hO�??�h��