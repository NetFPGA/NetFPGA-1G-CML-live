XlxV64EB    2b5f     c40<ĘJ~�3��=�D����b�1���Sp����H4eBxb�}��d��>ҙ"�.����d��tJ����+S"��i�L�*��I�&���O�@�wvU6�'b�ӑ��8�Adv2Z�,�d\s�8�M�k��8Js�2 �J*�JC<u��9�(l�"���_l��c�X�����(�=D¨AY�W +x��דh�:��b�P��6��5P��t*��-ݴ
6���r��_y��g��=��M���u_R��B`�ؤ}��o�]@��UJ�L<����4�{~�z�qCc�|}Q�\��?�e�?˞x���J��/���g����d5e�T�{����8ޱg��$�J��wK�w+�AC�ù�	�H{hA�/a�0����)�@�U�*�w��=.!���k��5>�p(~��zW�ý)H#2U<��cu���m)�ġ����C��'. ƹ8��8{r����8R��������~J?�g�����)�USQ-��+`H��\���Z�I�B^Q�q^��#���L$B���\��3��iN���%��F�����pC,��q�#�<��O���i o0`(j�Z�_zW��2J~��.q�����2��3x��t8#۶������ )A�mK5V��LN�by��(Ь����@8�.�s1���\@jN�.�eʹ������o@BO����nP��Y��O���x��O$��D\�*>+����@�B󲻉؞8[���pC��ހ��M^����M�
��#����r!���6T��~��;�<O��/b�ݗ�#��NY��G�B׮u[�����߸|���<����+}Y�ڞF��_ó#�3��s5i*�3Y}ri�,u
����ؓ����s5��Yqr�<�w���[S�r��H>�7�F���wQ�7ϰ+���+;J�!t�~�A���U#(�F��/0�H��tl����ר�jkPS���������t��V�U���͜��b9�~�!�I[U��/��B�7�N�p��vյ���}�����K��e���8P-г�wh����}�Q���|T/��wao@�ށ}��9F0A5qfrz�3P���*6��{���,,BP������B5��BW^����hg�Q��-�QN�� �rT�ˢ��s���&�ܷ|mޅ���(���~=ߜ�,Qa������pP$h!�IN��kL'�p����'�2+r�����{y��M;=�:���N*؅(�0#(�)/�N�<Y�F�јԵ �n����k1)X��O�/:A"�oG�k��>Ӌr �7��4�)E��\K�;�zOâ�O��zr����/��3�{Nxc��}�?��P��M��ٝS��������w�Q�~ap�Q�5��.�k+
��0c��0�����4�X�Ok�<	CPݯ.�vWA�&�'M����N��"��)��Ŭx.�W����e��[O���'�	'�L<ܞ�bm��yܶ��u�n'_F��������W���r�v����7�0�%��ұ��ZU�+@�.�Gu����gP�`��!��0�Q�5��@Г���dA�w!~hҲE栢������WL�I4�"�rnsm�G�u�'4��iX���\X�h��E�x��&`��-�3�߾��6B{��J��FaT��d�_+�l=?���p��y�;ŵJȫ��+tu����K�i�Q��(` �O���_hY8�������BJ�.���25P��{F���s]�X&z�V����C��g�A)g�7U�?7GpĖ7pk�~Ő4�,ܟ�n���Ms=�v��}�l�B��`�su~��j������j9s�-�Ю�W�YX��Ï�&��'�C���e yW2���o<�1���*�M��eKIL�7DM�SS�G�ۍy׵�J���:�o�B���9�v����]�k#q�t�Q�����-�Ď���)[���}M> �C��}퉪眼��@�M����ÿ4�ѵ���c\AF=�=}3̡:�ՂB�+�m�Cx�8\}���X��ś�'�K
7��hʹ��hI���6B��r,<u�$� �^퉓��R^�S�� �VB�ީZԢ���^��n����p|�#�Uk�K��8�*�b}� �'F��8"���4(���Sim����'WDß��E7��bT��BLG�RGc|%)��ѫU�M�M;�ҽ�����&�pD)�iH߭:E�V����8��_M���=��3�
RUe"�u-9��Aj�ߑS�>+���@�բ^8�N�/ ����x5=(�Ua���g��C,R���N�(��ނ�C�}M:����2��(A�4�­��XU�&ؽX�{>x��G�Q�6*��F�3���?�ycQ��0�4r@۽h�V�3�5���� ��B��/x��ش��T����5y'�?����g2�I;�=v�T`<C*�x'�%-���ߧ�;X|_1�L��#�HUc:�8l%e�9,kQ��7�ݼ���z�y�g�g�\ɿ���iY��%���[C��5K���ܻ&:U7�O�M��/�k�4�m�?("���k���-�3��N��	.!�Q�,���:Ի�������2� �ɾ۲U�c<�НX�٫����+���?u���6�:�-�㰁F��A���Z�Y�r;��%<���G���VAd�.�
6���ڃ?��G��@I��(-�&/z���A������K�Ŏ�k�# ���@Pq��4��4���P;Րʀk $���1��.\KM�]}D�CB
��h7}���tYS�ق�ȩ"cB��W�/W�������Ό�}x������L7j�]����ȋ��f�!���I�Ctt=)���{��ŀ��ZV�AC�n�b��_	F�Y����}>/uƻ�Ǒ��P�ʦk�����DI�Mʔ��x8�y9���������1P�w��g�(PO��qȈǻ|v��&��|���J��?iT��h���?�~��(�D��v: �
�=&{z�?��6������-&gr�����L��fi��sFYpT��-
�FWI���<3=B�f��}չP�6C�{���l�����e��U��N���㏪v��GG�=�N!{`{K4)E