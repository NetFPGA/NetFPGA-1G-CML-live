XlxV64EB    b8b2    2370���(���(8ZY�Зv�㑳��F�8�ay���amI�
�|����a���
j{4.�˛W�҄p�~���w�@S~���Ez0	�&��y�O��|h�}!W��hX�� ,�� s[]}�2�خ��Ng0n2��R��].���wL+8���$t�� 6��r6�o��4J��w?��$� �u���)�2'虶*zٵ������)\: Yp�_�����Q�(h@a	�l$A�I_�'^����*�rmᓋ� ��N�Va���b�,l;���]� c��|���D��G����Щ�X�^��_��`����b��ّ��k��8��\��CѧG� Cn2*�u	������s��A0:)�W?��=����C�i�I�Z�z�]JZ��Zk6�2Z{��B0�d��,�k$��W߁B�+^�AU�*WvY}׾���/yh�bD]|�w�a?���~������:y/�,/o�G}��b���WM�[x����|����d$�\��y��r�e2LQ�s$�J���C�?�^M�Ǆeڄ\N�!�Sn���0�i|�k_�n1P������V����(�Ԗր���� /�YVw�� ��˷@�8P�C,V��N�H�$Zj`ޯN���7�wa��>�"�0��ή����t���r¸�\�O�8͙L����ɯJ�×��z���gBāed3/X�qVy��b4�r$IR�Q���;��h����ղ�8��~��{EN�G7jj��Sм?�J(o<TLѢl��o�V��J��҄)���-hܑ<�AA���)m�q��(�X����a]��\�-A��H��Z��n7r&C.+�i����]�
��L�9*dN¢�9�F��:���67�zU<L0������Xd�-gI�#�d���f���>w,���n�A}�0�(��M����%����s!k�P�mE�h2I�@����>:¢s������Ht�|������'yܭ]ϭ�U�Z6�U��`ٔ���ȷޱ�,���J����N�3J4�>�l����@:컮�EU	۱;/���gwsX�� �{�[I�+�԰0	&��������\P2�#�l��Okio�#����	ق�+5t�y�*���am��ٳ���UsZ]�+Ό�Q�'���A�.��K�4\_�z���^	��)�{�<-��9
�Sm8��$_q�WM���j=�Qk�u
%4B*��[z�ͭ��1� z�+��ÔUP_q�3��!]z�/�U���$zk�?�[��c3{vN��q���:q�kk�#���MV:�.
&B��i1����A@1�{��:]z�jW7���������<DYN]� �3���kY��}_���l�˨<��k���]Z�ޛ�_i�A!'5Z�����T�
�ߋ��^��6�i�9Å���A��%�h��uyPA��݊$Ο��njőj�x�����qJ+��Aq�p?q�T���!�l�c�V�F��F��11�{,��K���d ���@<���u�ȯ9�վ�10�w� /���5���;����a�ꑐ)��	�>�ܕ~;n7w$0F�>uZi܂�9�
\iʻT$;n杖WeE�o�#<�}6����9����w�_Y@�_��p=o��Ы��]�٨�;�����z� /"�������E�r����{r����4� ޲����O-��鄬��m��nS@�6Kzئ�3��]3X�̳��,��K�]��oq�E�f�.�j��Ֆ{�q�kА�$��e�����=�!����h#�z4��h���Ip���TF_�݄�h~Q�&�V
�T�:�n5ݰs#G��X0*��W�f1�QcR<�ũ@
�N�2�����h(�ZVő7����iB��e	~�]�1Tp.Bd�>��/�B�"#�����#��;RIJ� \��6xW�u�w�.U��>Y���
K���K�x��z,�.�Yҡ/��\�Uo���؜��lۘ����mn�A�+�!nC�4��z����y~�`�~M��F�tRi&�'�l;�v�>�����ͳh$�����nSA�ts�.aM�Kaz�ф��2�����d���A=ʛ�o�TL_��#�
����!�?8#J:�t!t,!'�������e�y����udX�+}��wz��2�ձ���a�f��W��s耘e�X�&�f���<jT���Uݪ��kI��1>�dz��X���V	�'wꄚ�-�iߒ\^�GT���}pe^�@��l�U�L�$->�(G�N�-!�y3���;Do���N�Aۦ 5��\}�z����oV��"{iT�V��i��l=�e�E֤��-��y��H�[�!�ám.�)��{10ߜts��W/D�i�	���iM����G'�"�8N��fD�z��gW˹F�v$3~)���-K�;�-�r���s�w8-�O���RV!����tL�c�� ��%�5b��#�[��������cӘϔ,C��7�$HU��fRz�F"�77*b��e(�V��,V!��f_��$�N��x�& ��H��������b���I��}q�҅ڥ'����/&���8n ���ڎ�<&=_��d�����#m�ڲQ���:�3U�A��pͿ	E�Lh""�ĦY�.��}�wr��^�R�M<��V1�hK1LYP�U�?L��^�	��0 �0@eCn�,3�$4�si���E"W�dX|R�������SJ=�$bv���/g��_���g0�&�k.��S���'A�FFyS�W��Q5ۨJb�tqO�)����Ǿ7�B`r���^�W��W��^�����/+���d��%����>XԱ2��CU���]�2��
��B}����x_B�������a*�<�q�6����7��G��|�7�!ٞ�g`Q
��dh6��ϸc�yr�#��*�HA�â�DmǸEv" ��h�I�(�<����V-/��yL��lY�!e��E�r��s��k �b~��u�����a���l�&皤wl���̖�I���ܱ����"�S��4��S��懾��p����c:N�G<��wĵ�x"�1*�2�������n���U��d�Z���ØSYf��tڪ���`NF!1� )/��}5�$m���3���o��(j��vF_���]$���}����q!��-z�<���a^�tU9��Y�P��+e���g5��I���=B+6f�0�o�f�O��ͻ{L��%D�{
'qi���=9�|��2:0�_ّۧL����Ÿ��f4�n���Af���wf4�y�>N�j�Hs
�̑w���� �W����
��t>}������Hq�,<r��7"�u�>�ܵ�_��$o����Fr����Ėr%���"G�|�(Vkb��q��_�F�^�V�N���W��A���TNr�vqa��Y,B^��g��Ó�~I��c� �Y�g���9W�"M,Ո?�.m��ku½$�c��I��Wv��H屒>xϓ�f�DQ�N{��@�y���5Қ,t���m݇k���P�L�M�ݞ����V�b>��N'���l��J�Q>|ni����ty�`
_CD�0e�t��X������3�ɠy4�5z��J�`Fy��N�R�����c�TS�K��k�7MDE��@JT������̒|���"��e������Q�oՈ�r[?��ݿ��=H/�I�� �S#�v�"{����aC��^��Ӈ��֝�t�#�v�. ����`Ď)��@��`�/�i�H��rl�=}��HX�7W� �!���=���g]Q�;q73�7��I�L�,�Ö��Q	J���{XG�؛�)��� ������d�A<���g�@�_���\;T�%}E��A�@�њYqT<tfN��}13��߃�bdI�D����`x�\�D}Q��"������-٪��T}$Oc��u:���O�C��ow�G�ر�9�]$uq�<�}�*�g�)���F1�W ��=u�3Į+UZ'<&^��Y콢]6V��>�1�L����>�`Y�G�g3��,�Cv�-)�Pfc�J��];l���U����r��-.!gA�!]"��,4�d�ʥ&
���ox����q;�t�NG�������)���wK���5x~�@$���u�|P��a����e�����D���&^���"X�Ӳ^wu���aqٸ�b���uE?�i,����f*�+���F9n����^n�[�V��,��>T0s}(M�gm�~����\Dȏ�ь ���|$]�X_"��f�$D�{MD	|�]ɖ��z��������3�xh�"�Y6��N)�<
�{�hW�
0���{4����|�E���%�TzV��K���}O�POHf<BWj��H¶y���o�g�۷���2�ß-z>�Py�nI]��X)H��.S�8��Z-V�%���&E2��W�o��x"��	j	֪.ϓ`�ɼ�r�|E���E�Y�+߻G������Dss�,M:)���;��__�:����k~=��yiz�;��f#{K�L׸o�-���s�T�Mx-054�zj�ЎKS��d��x7��9�~����2�&u?>	z�B5���C�m� �Ҍ�*/�^��F�䑟)㝥�������0oOM0(�dQ�RI��J�	v�2����v䋲D�D/T�Q��j����?im��&�j%ذ�H�/�I�5xS^��r�'-���+�
��n��S��:�+�yb����DXt6�B6�n��a��UF~9����jd	G �[���R%B��M�㶽p�$v^�,�����!��_��t�:�F�M��tG���S��hm�N��Od[ȫ���n��ޛ)"�m�������
��ےݻ?�G����0�H�o���A��O�R�7��ʬ��<v�iבU���n���f�����,�?𗥹ٷ�'h;p�~v;쏑�d����Բ7pB=� ��%� ����Nx�R�)<��N|����j#�S٤�;���o�)��lΨ����|�d�m�͑���#�Q@s�|�`��7ƨ���}",�|�Sk71�������㊅;&����m�AgH���~7�R����6��&�Q n<֚Zì��zr�s�M0��a���mG0���q%�w�dv�=0eg��%:9;�iM��փ)����"pf�~3���w"95�o4���E���r�P��A$�'��<#������h�(y� ��R�������g�p��'e9�}�޹wˎ)�qEofP�%K�A�$5���la�E̱t�I�@'܈n���t�JH7�%AݞV���h���7 )�%p���X�v���̮��C��e2���1ɚ̺)h�<),��� �w}�@%od����1VU�rl���
�_���K+U
-!��
 -�I_p���ήaai�µ�*�P7�V2��yp�����8ql!��ۉ�b�.�ޫ�j�cӪdZV�#O���z�a#�W4pkn�.2�M
�����pB;$8(�����8(�mv4VQ����L���p�v�=�1�EkJ )b�!3�,U���@)�ܣ�����y������Ť�'�8�����W���V61����R6d2X���]i\}�b��*�+G�"���b���{{-+��x�7%�0K�v��a�!\eW���D����v�6p�b�-�'�\�<���;�J�k��&Ҍr����j1�ī ��3$[�[�W��U����;>|�t�翑_�
}���D��S1;K2�8*<N��R�."m	������h��X�\��&�xK��&x�N������dX�R����AO�A��g�r��P򛇿����hj-z�y,ӱ\Щ��S`۲�o|����΍=��K��*�?f���Y5--�1��,��̞�����%̣Cw^��3s/ɔ f���9��&od��i��f4�r>Iؿ(��ՙ������JS2=�*Z�����dXS��l)A
�� �Z��d�������$�ʏ�����.rzRS�q)�:�?�6�؄#ݮ�6�����j'�Ý�4K/(F��o�IE�[��~uFF�9��#�ړI���z�J�8��o���#ӷY�ak��T�;]��`���S�Յ��$L>v���$�0�z;hf����8�w�Ԃ9��3��a��8V���H3v����Y��c#(�=��6���k���fԅ��V�#Y�I��n�q��̲��^�&!p�����Z�6���S���<�}Db�ABW�/r��w[�m$���a�}�iC���j�f=����i<���l��qTl���Zak����{j��M�F�f�}n�S.�ittG|n}ZxH X؞�%c���s����JO���FīTj�Iw�wjB�&�G��,=��H�����`
tې�)�S�g�г�N�c#%[�єj1�<�E>���l�h��z���<�Z�4�Zȟ;
M��1�V%�\2�JO�\!�ٶ&J2�M��Ԇr�CW�����.�8��u� ���T����-)IP����~ik��+�ȩ�@R�;2\e|)��QBI�Ѝ���Aw��0|�~�e1�b�2�̷ɛe�׻F���X����H��꽭 rԈ�ڟ���~���vL ;�R�WRzy;�{M}NE2�O�[x�2gt6�q�:�>A�YJ���]BF����O��@���}D�6�M.d���Ћ��?sӡ��D���r�R@��]S�M�^�av���'�d�؈K�_P8���'�`.ӫ§q+�cڬ7I�LK�����.@54�o���䒜mCnC/�Ԍ%'�n߅��*s���YwK�=9ww�����L��6��֕7_fŬ$f����Z�bJ.B�������]3jc�pk���~I������B�X�U*���X ��"����TЬ��a�|�k�_�0��͵�,��B{�h����\G\�R�$���,�ܬ��X?�rrTWR�����`c��#�aZ����m�<�&'Y��t
Ę*����Q�XL�f����A�O2H����ȹ1U�A\��	$ ��I���%E{� <��˴�Lw]�1Hk���Am��,��X�̗ �.a[��؍@�������|T�'����_��&<�(�v���e<i�a���KBTj���o���O���u���Ns��?�c/c��/����T�!!e$ƌ"�L��W�n����dJa��]�Sw�!�(<�b�֋$�p����EL��2d��49��{r�#�VMO�
�sˡ2�1�H>� �����'Kig�	} ��U�r�r�B�b���C�������A��\CH9t@��e~��s{��Y��.p*�z�ˁ���l�'�����P�B�-|-ki ׊Zĕ�S�+b��wեe�A{�D�����v�����if��{:O��:Z���T+�����W�����jrq.�L�"��O
i�Z	<�+��P(�Gn<�n��F?߼"I�W.���s�d�-�,���6���D9����l�o~��\�gP 0��"��?�� ��k|W�΋�#g���>��^}�kf.����d8}F�DQB�J2�Y��Mj\��'��ﯳV�s�N�r�=6�5X�[(�݋@ 3���6��u��`�6���J ŹI�6�!�L��Y�a1��)���������U�̒4��}�*dѰ�_���P<�L9��7�֝��JR���C�&�ܝ��o��N�"���y?�+��}Ao��sMD�	g&�.i��v�����o]���H�ڄ�H�jʗJ���v� �0��o�����T��x��[C�X�!c4�_� /�Nm��+؞>��w|S����Y��T��K�� �m���&x��4��4���<j����wB���N�#n]Px�S'kv,��0�g�f����|\��%&�仨OA!�v�jN{�%I�D�I�f�Z�̾�jqB�+m�������T��l<��Wʷ���U���|Z|y���$�}�G��_�; _� >�� ���H"�Mq�=Mj�zY}�����7�i�.uL�5�/m��ek�y�����&~����耟��*��V+'{x!�'QTq�#jA�Dk�2�SM%�3�I�j�>�8�PE�z��$�*|8�/��Pĭtn޹�Q�.S���Io!̧���P���n[��	�,�"�C���_��ID�0vhg�ʁ<t��g�t�\���Kr��� �01ۘ�E&�����I�`����V�<Z3m���϶�䜢k_�x(�(600*4�{0	(dY1���Rs�DxD�y�SJ4x)��`i���s}��!��"���g��a�J�F�B�_&z����#�����]���N��tBY�~�)�]��N�!��A�r�Zy��rD�
�cu���d��S�#��
q����$2�=�2hK��sd_�;p�
S���u,��;i䬬��
���5}�J��W��ށn���&�l�VJ�y��T�	F��T6��t���A��_kO;��;O�T�֤b������ RT�=WҾ�J�X��( ����G�E!A�-��m�� ��"�s�%�m\����qR����d�j�7p}(��ۭk I��d�)p�=?��x�8`�����T+�
�w����;�[A+��g=�H��^o�@��o8r%^�%�}�30�e1�J��y�EC |��k�Ds��BsX!W�#��5΁i4�J|_�_�_�͠��zhpk�|��J���v����V<Q:b������Z����%��� �;8�y~�g����&��a<1m�M3h�@��v�?ޗyg������W-��Ȑ���<�ٛ�*r��jd�s����eG�S��{�r����<Y����Y_Y=i�T�#�I<����Ӛ[0 