XlxV64EB    472d    1250�4d��`�㾝�(�B%Q�-}�n�m�Q����9+d;��������r@oy+VeBn���b�`.T*i֟�,%h�xl�8�X���G';�J��\~.(�������ۏ���mQ�/d2��@q�Lɩ����z�e���*$�D�;��<��j����y3�����r��]?3�}���8�O\��|<��8K��� !���D/�S�4�!c���������u�BןJ����D�A���?a�o��3��wZ�)�RC��^@͛ҶOa��j,�bg=M����y��$њh�0R�T�y��پ:�n	����Vg���Q�ҽ�^�\u.�f�}� -�1��J2��H�p2����T�g{M��e`+~�(���4Vu�V��&����Ő��	�_˫�@�ѡ� ;چ�f4�~��K�ڢ�� ��T��u�T� �\1�]�o#&�,���Dg�Z5�f}z܋n��*£ �߳6]A��2�Y{pj�Z�M���������,D@�m��ٜ���Ɨ|��{,��C�+��,�+���=T_��lz�IH�9�J�� C�O���\l�+���v��I�/��	�.jzDo��u���[1�m�/�
��O�[�R�7>~)
R ֤��za�M����?�y�&K��sw���4�A��T;�����A�����,'�sCJ�T����՟6�i�_�S�L��H�?`H�I�l��u��D��k�Ibm�gm�Wl���m�����%CI��-\M`���έc�M�Wj
�5pt;r������m����N�\=Y�"���x�r�NȳX)�Q�����G̯q������hFQ�Y{�H+g71���]���wd�&"��y *u�N8�8*���7�"�cx�2^�ɡ�k|C�*7�F[��r�O��u�yіo����{T�	˟��`%����rT��d���;r3�#�Jm@��gLXU-|� ~�0Jb`�1���J�����L/�x~�X��+��ph�~)��	AS���R�J���8'�u�#�UF3j�2�oy8�䠖^� ���lc��U~���X��D����:��P���6r�c�HP��cO&uʮC)\�[����lЏ<b���x#,/�pfB@Px6���f���2�T)ŬX�s�B ���嬊{����>,�ņ&��N����$�=��J����~�ʡnJk���u�����>Afwe	�����4h���U
n.�U?:�]����?�@��oq{۠rr��k�;U����sv�P�*6׏���2t��w?�����M�h�/���][�w�l� L���ޕ���sS�C����9	�N��������.$K�(=��+�!qÌ�.�m1�y@��KK5�p��_*���N��D.�y����v��O��0�/���3��{B5eĿ_��d�|<�*җ��?�i��.J�+�����h>.U���K�d���h�-FP���V�:��dܞ���ao����Q���/3=�.i9�%��5v��_�3�+�	�����;͓M����Awb���
x�S�A���H�*Ki0�x{��;-��ͫ��Hz���^��� �pnW���x��|�~�����9b�,l6�Gfm���A���d�2{Fǔ��$Ҹ�r��9���EJ�EX!IT���d[:L�-l@���qŞՎ�U��w�ҵ4�<S�R܆�eQx���>��|���$��qS��
B�!�߱P�h6e�.�)��UL?tX���s�~=���5C����>q���qk�X�L����"˔3��>�"Bc�I�DC-�s�
�Cbn���WA|�е��E��
���N/T����$���r)B(C�h���Ӡ�S4�4���Ԡ��/��}��L������������D��_�ks�DM�����m_7Q��*��s�N�����_!���A>�c�Z=�{Um�P��,,(,j�W�$��3���y��p�`E��|G�fxM���� cCUw%+yC��0�e�U+�s�M)
hv�Ý�>��@��k�Xv'��e�Ws��*�d4p�̲ض�ݎ\����wP>d�����$mf�S���{M!7�r�-�7!�&���������K���zؤxe�%PHM��$ﴀ�R�P�}W1�=O1�u�s��'��r��
�{'(��/RS�AMQd+s.;�o�ǳ;��$�0Q��&���!4<\Z+�������T�;�m8�hB�
�&Z>u�g	��S�3[�y�G]u�y��?<�z��][#��n��n¬.�ɶ獺;�� d���zם��od�͕�!���7c(D�D�Ya�z���c���8V_���c�n$���.�P�~���)��@~���d�U�=�i^Y:/y:�$n�E �
�3��~(*?�L=�/�_fh0�0�,�Kw~ �F.��E<U�t����V��/�蹣K�Ce��.	�Zyo퓢�Y2�z�pP��'�Fs��}��~s��N|W��;��螿��R��z����M�������G&�dNnL_�k�R-�8�L1�O��w��v��בhMFE��y���s�Ÿ31�z{|_:�t��̔>�Y)vC��z�����J�ٽ%}��;�~ k(���K)	P~o�*� �q�F������2_��c��SYƮ9:�T� [J��#�(د�7����SɿKV��x�׵�����4�Hډ+�~bw���Nݔ�f�H��	�~�`"�v�3Ē�f�5$�U�_M���X��jQ��z�Y~�� j�L�i�1SQ\�����h��U��GD�k�u`��mE�!<U%�hV:�������ad�-�]є�K\TL?���(Nq�#�~��:L��Cl/
 �C� ;��~Mo�-~����g��7y���ʌ��\�"���xs�)�t)�dh���r��Wj-��^�|-�v��Ke{���i���J�䄴�rQ��d�s�ve��Mwz�Й)�񁌝ԯW������U��z���R��5�)��F�ɶ+{�(ɠ��m�6���H��y��vj@`^ù(7\����_���b���q��[�v�  ��8��hO�J/N=ii�l|4VR�n�xWq`��հ���mR�"�d��B�a�9,����Hd���6�ãY:�V�3����D�K�ݍ��������̩B���, ���K��g�V���,1�R7y���V����֡,�m^fi�H̗?�>���;���N�����J�$��A%�(��6�hp���"S�1�M\nK2���H�V]�wv�*uR�׹�*/�������W� g����o^E?��)�'LL���쏡N�E��:4��.Jxug�B~�LfG�i��]���9ɐ�P�یOhu5��Mҁ����z�!�������@�q>�$\��Ǿ�;�m\�f���Y�$��݅�8���j
A��.i����QH��h!�|!r�8���瘌2���1�.�㩯J��� ���%���+�P/��4`�hL����j���,�5��D��Ms:F <�P���|�kS���F�?�N|�,Sf��i����{�"�UpXF�gͬ� �,'D?+���.h���:����cTw��Z�z'��p�S����0H�9��jk��x3�����K�pD��ϻ���j�F���c[������ɿ����G8� l�@�{k�.\9S�s��W��~�GO��!�l|��ce\E��W��fJ�m�;�W)��G���Sn��ɕ>���?����V�4�Ѯ�c�_Е�C�Q=P��[�� �j*�?}g�a��J*�f,���EL��%�1�U��t�A��[5�i�\���䂘b�1�{�W姨}٤<�)W7i��D��u)B�\�0��̌�٥ݿ�Cy���&��n
Ğ��h�����痴l0*^! �(t"�lf�l�L�j =Ai	�!8�TU���O�笵n�|u�qbr(�;KbEvS���.��byk^��D�����U�� Z�p���\'�R5���>�|��Y. �(��|��T�����x��61Av��(�>X�xʎ�D���W�sj�����p�)����o�_���coϼ���/��J���è�wi�b2��τo1�pt1Wv�+�Ŕ�oO�������G&t�x�����M��,ӺT�Z���<˾��JbN��|�x8�Is6�J,��*Q��K��1������� ��y���^/н�Ӥ�\�4Xt����;�į�%�������b��G �����,y}x���c�B��;@%��I��܅�B\��=k7K��n�+�R䯁�V�>��+�CA@ަ�\c�TFp
m�:�t���|��Gy�u�5��y<7�QدJx�_KiO'��sq�Kf;qt7ƛ��K���A��M��N������쮦���,~�oq��*�_I9a�Z��Q��ؓu���ɵ��Np�L�l���H.7�-�]e�	s���+"��v��d<2�OҬ"	<��7O`7��˭�,�8�y������=B!�V��,P���F�.oO�\�RܺV�%�/��Z�y�5~�.[6�0��S�!���f������6��@�SԸa�(;