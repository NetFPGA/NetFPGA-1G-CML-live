XlxV64EB    62a0    1710�=�ǊF��,���o-�n�M��g�{���[��^��h�G�7���xWu�-q6kS�t��NxSuƯߚ���TM��|��ʢR	܎��Ժ�v��3�JU���G���	�(��u����ŰD��n<P��{�	�r%H��e<�s8#��u:�2G���d���s2+���w���%4H���"ry ��:EV�_�D2k��y�����T�k���7KZY�N_�O�-i��v����=�Ĵn-鱩�b���b>R�H���A��*��]`bǾs�[�Bf"���5ݗE��dƾ\f������d�[J�2�p��YY)$��"�72�i��#ڜ�;��ǩn�cj'm��.��S��p+n*�L��%O��1]@qv]UX*Eg:V�ıRL_�F?-��ȝ�M*�+9@�e�p�����2�$#����Z௢���.z8�8�F����>z+2#1��Qv�i��~;�&��@Fi����)If��0��`*!?�����Z��|ҵ�:��E`�$4�s�9	2��w�pj��xi���)h}N��&� r��l8�s*|���E�	��?�T��=��G�9�)�-�g�=�X�v�D�=���(�h$y6��������1W�NC���#B�͘Y7���	�� ����BgAC�0�����\3poǲn�%.�c��"\�l7�7>{1g􆳶�wښiڦ�H�S� a�9���'>g�9�e��n|?},5qFP_�\����Ư<�L��YTd�^Լe���tٹ��d"NN�W}zP(̶[��h����x�>A��N}E�	"h�^��
�;b�9����?5�Y�/WB�H����CF���X���d����f]�@i.d�^FDn�xO�+pj�d).�I4{p=�����TY)��Ъ�W��0L��,`�z��gV��S�S�J�!X)S0��F��zJ��@عҸ����C��a��Wl|�6��=x� I:�ۛ��r:܌�ޱ�A�/i�jˮ0�)�N�����*����	��j]�2b�ޓ�q�<�˨|z*g�o�f��m�����ġG�{�A!��m0��\9O8R�OT���?�T��I�M�U���~�0��3�]���ǅ 7�Ӕ�#Ӗyƚ�����	�UL�q~eN_~��3H%�R�D�J6N�"����&�X��>tYД��}`��yL�V����!�=CZ�6ɮ[>(�U�@uJ�|�Zնus\@�D\TS�U��e����HQ"�z��	�J���YA�hj����H�:?O��NH�T2�-Q6:��1��e:-/6����� ���� @Tž�����o��XO�|���G����$x�t�d�i������ϣ2L�N�A���Z~X���Xŷ? E�U���o��Ty_����v��6ٞ�α��K��:z��ǶU�����2q��#Q��K��N�5d���W���"3�#�Cb�&�"8��P-�g���7`A(�i��<��=��v=F�l�uF�
�5�
O��Zf��B!Z���v�%̖F
�b��Y!�]���6X'����&�Q�� @����56e�[�n.i!��~��6<�b`d'V=0�&�D̞������ΊnżnE��|��tҤ�7>1ؾ��CIk��-����"�2���DK\��-�`K��5����I���2�d���y΋1�������P�vwj~MB�$�@'����t��R)(TD-�1��^ӛ��(ݕ�E{�"�T�s��
UNuU�!��j�p�w�Г4�2���Ca��N�j���L�t~�Sg�K�ʲ��:PȢSl�Y� ؽg�+��<,�J��c�;t!����W�/��Ă����/����~v��-��'sv\d1z������]�`�ZXJ����_,u���	�����[8�3£LfwҜ�@���y^9H$��Gs����l�{�'���	�Ky
t�Dg7��N]�qgH�� ;{1��4��j�;�3eք�a��pQH��t�Nd�mP�(�I�����o38�Z;R��c��WU������|��ɩK;����7��n�+Е�O�V�捵��t�ڜ�C��qDA":��Mn�H���:�3�@j�L6S޺H�'F�4O.,@��`�
�P��w�Ԃ	"��;��,c�v��P�9M�)r�#�Br(H�����s���$�^Y���d2�u�4�������l->���z+��b�S�{��m�%�JLS����� 0��E0u�(���^���,��D����T�+��0�{�s9I�����a�"�a^7��փt(}�D��'B\��ۖ17=�����8k�b��b�'YG3W^��G�{�z�q��yl�}Ӫ#[�E'�1�蹼W�V������d������|X�����r^!�2G�"�}h�S�Q�u�k
�{x��o�m2G��|��*K��9�ER�¾B��ք�qޫ^n8D�P�}<�9�Sw�6�6���+zXgA��g���z	@7`�3F'��oc_��4`t=��0cna��ַ���F�7�qB�.ߞ4��.LO���B��@�������Z1��|p�Ud�'>�vpb��Ï(%�ҹt��a /ДG��k{��\Gs �λ��N�n�1�ȗ
����7�����x�`DK�زD\i�>���-�d���:cS\��7����G>�ݟ��\?!�����uC�XT7X+����0[�G��g��J��$�q��3թ�sF�d���@Ap�JL�޶����9(���!�m�, ����Jt�y�aIu*tz�j��onB�:��g�t9����}ŋ�v�t_�U�x��R�9���G{�6���b�����2��{j�W�j�x�2Fc�mw�q��Q���FHZ���Q�մL2\7�����yj�	4�Gm�V%xr���n�K��t��;%ٌh
t<�Eۚ���(p��5p���4R��0cj��:tZ4JZ%$]�!�2-y�r��~��{P~j��һ
��b��Ih@�/�#tjA�|9(�e�wSx�����g\�
w%Ͻ\������B�0e��J��*P�6����� ��+c�8\e�ud���9ע��8�)��	�ԛ�t��9�5=�a�.�g���uv&�!R�&�*�q׼� K�bV�Iձ���"�:���}�B� ��nt���h5���=l�(�4�
kT�zT}�=���=#{a�H��a���b'z}�N�~�%>��A�8IF>�X�v�b����B��^Ƥ.���@Br�N�G-,���_9J�HjGp�R?���tW��f�1��>�GN:#��������	�$¬9`��q�},j_��a�Y�pZ�lq�l��t��)	�V�o���_ի�^/f4��
�ց4H��3 �S�4苈h���a���������r]�������r\�"�!cQ���ȷ%��)il�/Z��4��8�(�[`/2�S� @���+�Z�x���s?����X��G�h��̓)�ϲ����y��:���|��,�+��^�6�fPp)#�����R���}^���(���H} {���'�]:"v�l�#]����L �:�$E�����ũ�@�ފ3&O锡q�E��;\`J�Wa94���ڍ���J��ǿ�c��\e<'�w��.\�a�e�#�cSe9�e��fr6���]�'��c9�XS���H�H���h��1"�S)��e�c�g�O�5��\���>C�g��r�������u7�����F�r�/��oSz���0$���௙�N�G���Y>d5\]L���W'<+a����Dacv���F��'�d��<\� ꘝwo�ܣ3�>�@t\�muw.��-����[�?�pb��{'��JپV��$�w�K�2=U�m��O�C�(�%����E�|���]"�)"#�`�3z�-7X�P���|V^̬?�0��gR��?�hc<�-����Oi�9A�1���c����ڎȫ�x��B��v�E�Hg�k�����s��ERk��s8��Y��a��2���z(�oE��Q�g����i3�3�dI ���s�� ��� ���D&�R"0R��"y�݂�LKe��?�,9��ʂ��������o(�E8]�'�T�)-Q�d)I�b���]�n����%�;q����Ӹ]Ya_�Y,�}����sV�m�_�:_\B��(<rVz���s�c�6�&�	X��t�qIQ�T�*k0�钩*���҇h.����"{_�r�W�H���v<��&t�f�K����q^��J�]�'������-�,��+�ĩ��1Hb� ����uɢsib����$9��^�2�wҸ[zF�r�&����nT�2�+ó�J��
���ddt�qm�5����} /�`�>��_A�of��ˇ�L�?������..!����Txqd��qn
��_G�z��4'K�7􌨣�B<u�;�?� ���]\\�1\i�������}���+o����B��Ͽ��I��,�5P~�/��uW�|f�[�����[#�.0��X�-���K��\ɺ��@�צ��=�7��SA��荳�HGp	0l��>?p�~^qi�0=0l'�b�n+c�hⲽ*�cK.�9�0ny�3~F�1ז�R� $9˦�o���vm��"�qK�J�0Y�p��ڪ��Cy���i<!#3����] ��!��#-{����ZF�A�OZډ���1rE��2�dٻ���m]�ڨ��Q�?l�;��h��9J�T������.���a(��L�l�]*x��е�CFG)vL���`.��Knj����"T��p#�k@R�k��Z����`�����bo�`��oG�O1^��4ܲ�D�Fa�;1��)5?d���t�|3�Q��'h�-���s��Z�"0Y���5����U�Ei��Psfj^�߾����gN}��9e�3	-�l3BQ�RyG��0��:���:�|��&b�4%x�������aS��-0�(R�ߛ�B�U�z���x�#�@�-���y}��,Q�uǒ�C�������H�6ؖ!��>b��#�g:t��^A	���e�f��ԁ85J���+������2n��F�Թ[��oi��<�l�s�$ܦ}?�A���#h��9=���j�L�4��⸜Le��6���L֐�we.��10GZvI<5v��5�D_�� �?��:R�������Ӧ��+V)�2���f �������R��?0v2z�Mb�X� y�+׫	��z�H1c��t����6s0@���������+�Y�BV�3���L�����+M�QSZ�ψV��c��X�������	��_K���y��O����<���74��%�0+�����ī�X��L��䗠hr�w�ݱe	W���r��-������c�{|
�E����Ӿ赓��t?VF�rϕ���|�>��^��u+D��po�{��vˉ�6L���Ԍ���P,gHR���?�V}����z̵G>W��
kC�(&�f��X!��X��f=(u��ۧi�n`�C @�Ab�QT�k\��0'#��r�˺�y���Ɛ�j&�P�'�I:44!~�r��^b������^�z�'������""Ωo��N_CM�l%֓O�S�$���Yi��:b*NIf[���o�yy�N�n���T�m$!�$b[Eo���?Vr�q�V�/�u�Te�Dz$��,Kf
�z��/��t�W_�����FC�0�,�A9?w��`�/�2�k��Җ�������P�Lw�]F�OM�1�؅����o�(]\|�Q�