XlxV64EB    55ce    13c0T�47��ڿ������D`J�Ѷ~�NwBeo��$�t���M,�xM�j�r�"�5�;s��.�?��Y�o�J�V%�� ���gJ\���woT� BUK��ۈ����=��*}��,kE0aX�vc����B��d��Gp�9a|J �?���*��X�AC j�(a>p�i(&޽�6�����=��?D]���.���"����L$���}vO�fٌ�z=.�
 ���Y�A�!_66R*44�e&��1�����*ha�{�]m�3�5�����yÈ@	S�4L��	Uϊ�bt���c/z
}�	Q�
��_�Q!�H���tQ��Z�4*VV�Z⿒�1�Q�~l~ZTu��M�C�Q-3�-)2Ȕh��䦌�Ԑ�_ L��Kj���l
�%����'�	��b�����"$����k����q�������} 7U�w��'�{|���7�V0YD��g�KTG_�f�a{��	���#R�Į����JU�����M��	�o���)�z ���E��8ذ~�R8�R���������)y�Mf&���Cn��Ŏ��=�
g��G�ߦ��z��!�n��2(���E�Lb%�~_T���L���&e��ń�z�pI� ���:Yط�=j+]Z~�i4$�N�����>�qӘ(��beo���,���d깣q_]�v�ԘWz+}�:G?Kɏd�����^+� ��uw��N|/��Q�t�A�>#K����tc�ym�iah�`9�e ����:JW&n�F�j��<h=20���rѯp�nf���P��d�9z!�S0!���	�p`r��6�G��hm�Z%
���L�M|i���h�.x����X����<��F��P�!�	�gX��,��Uᒝܨ;��8Dg��Ƥg�m/YT�J#�����{E�;p��/�Zru�z�
_d�	J��ᠫe�k[��K=��Ŝz�4$7�FWv�|R�D2���9ì
T-r�N<dj��f�������C���G�a��ú8{v��W���o�O)ƨ>�{�r$!�aZ�Y�R��~;�7�Z޾�HMn5~|���.�+Pyk6�
��m}QJ?^?�n�W�Qf�`m����ljH�.�����X���O���[C��)_h��9#��K)4��e��0&��t>�օNɁ��/J�֠l���w,L��sh�R�#�7�9�Z������k���%�e����{��Q�;��ӐwaM�3Au�1u��ٮL͵#�<	cT��A�}�.U!j�"�2{[�"	�>�Ǜ���A[缼=�Mz�.������4�A�a!��͝grp��%�]�2��`k�@��"3�~W'�[�rc+HB����hK�P-�ꌤ��ht�r��c�X���b�#��3��#(��G})؉
�'���!-.�(ys��Cw����=B5.0�;���;��~�%��R&�dáh���TW��O��&�G7�Ȓ(��%��R1���5�<�@4jY3F��>��'����Q���02jx#k,�v��:)�%��i_��p�l���{C�ǐ�߰&hR)Yb<�t�D��/8�����s49˱�^�����r(�~���.���f��Y^i�v0ڑ�h.<p���
�;���>Y�~�Ux���bW�r���Ԍ�;��PY&�7����N�R	]!e���8�w˙œҒ�r$q�0o@#�^%/o���*}�4�Sy�U��WG�-/���Uo�GXg�}0�a��������޹a���v�ZP��
Mr��� c��#K���N��e�̘�hQ!9q�%̊�D[=��>}��?a]�%��]�U�{z�3+6�"g^�ȭ����GM�n�O���v/b�9�bErkh4Ƿ.������Yv*��	�j��[����4�=V�G��m�z�<�:Y>.1"�U���?[�yF��BE�Q�l��D���rfm)�"�`�2!@�ۭ�H� !���h��S=�8���cg��W��P��K�8L���{ŝ���$U���FV�����kas�J/��l�^M��H��x�ȿ�\��j!�P4-���k׾��~%,�[L���_�U�>��zS��"��a$���#�ΡVnU�"������:ي2|�4`�hw���3h~��7+���Ƈt:`e��I5-Cm`��ҡ_'zJQe��?���3?� Y�2���,d�LO�(j��@P���LĦ7��'ͦ|�q�Ǎ�J�~bƹ;]$�Qo���x@5\I�W��H���\��〒��&�Z�"`�:�0@s"v�ںZ�!'�^X��Ң4��/�����+��m����MJ��ذ[v��PIM��)?�q�34`?����� ��M8�,f�8�8=/��~��j/�&7o��
�N�z�.(�[f����?R�&�Ġ��5��ы��)�Z��<ڕ���b�����d7���g�t��}#I���8�'��T��J�2)Fh�D>�f���;h<��#*����0�0:���E�DmA�L���f۹1DO}���m��P���C�=�奛��VS�Yֳ�r��sф�~�J��ځ� ����*:���ގW�\�3wJ$]�O����	F����N��4�M��}��Þ]B�_7����BՊy�!�Yi�����ܤ}�P� �q.�@�)�n甩 98�LI��6��lc�*vP̏�b<Z�C�\�Ad���W��.>���J/�Y	�+aȿgE]u��K�~�~�[�g��8��H�(~w,�Z�;]�h�yJ�NiN��`�i[�Z���t���� 3Q�臄bup��+p1������K�O�{���d���pc�e��u1X�sm$|:�bM���x�ӷV:�:\���I�3�W�aR7>�0��- �<��j����"�q�8�@�W�X$^� W,#�*�����{����r9i��Q��Lcۏ����s��a�a���29��5�`L��f�l��U�䍴3Y�D���9�eQmN��~������Zs�'؉��RPs2� ��\;	�~�0�'#��ˎ� �J��oKx���_��_��<⪵#4���hs.W&O����Z�����վg��H�)
�0KC�yq*���T����U�-2�]yvʖI��LG՜y�H�ĭ")�1ؼ��o؝�XRWt�%�U��kk�QT��ڷ������i̿���,^�DQ^���B�8�"]%��3�9�������%������fߖZN�W�Y�u�vsh���pHZqBt0z�>��_��\D�@8{m��!�x�M�p���ti�	��y�^��N��jh�g�\k3�O��u ���Nl~H��0(e��(��ɬ��g8T�3�Pѣ7���#�G؋:V�\�����3�{O�ȋj*o��Q�3MmVJT#����|�Ս�� ��Ő8�7�$I�׵o��Q�ew�Q������2瞓
/�z3�Wu�:�w%`ś��+0-�7�	]��;��wb�|s�����.m����֠�����NV�E�?�v|^5L�m(`"���#Rҫj���������	H��r;y���]6��zg�(ݵ&S�(�{nR��$�� v`1$��U�My����\:(�=@�3nl8V�0�������bB)���d�<��I��5��H�Q}����ƙ��}�[=�.<���6ذ�|ː����*h�c�LM��^ʈ+[�yя�~Jszt���j��&�L�Z��"?�ώ�zs���5�S���H�}}y����FJ�G&rE�����4[��ח`�5/v��{ ������k��(Dq�?��Nk��(�B��^^�,u��W�D�I�ޘVV �o
*���fh��'��Ʒ�>uu�T����]u�Ψ��i���ꊏ8���:�� X(���ö_��c*��y�d�U���z;{;	 ���MF�=\Kya���,�)�
̓���,:_��{����Ӿ���B�|�%urU?�y���Y�9-Q7��?��Y�e4?����΍���Da���}>Q>|�I#���!��4�Up-X��Q�ծ��x#,L�N�̠)�#�@y.nD�Aq�k(#�˃�saICC�S�ߔ[S���YVt=KC�$*�0��٘�?I� �U~k�.r?ls�?��PA!q#����5[�یc�v�� >�r��+\��v�-Vy4��WӔ�[},c�ܐ�I�f8�j�2w�/����c2LO�ֿ�>���+�_o�%����J��� XB����u���-R	�Ic�QpQYޟ�9=�@�H��-�a&��Չ�<�Ӭ�v��
��۪�t�(J���@�BY:�{,��J�J�n�m�$}�_-�%�%�A�����@�ؽF�WZf$�#�F �Olew(����I8���ӟ�c��9�@u��8�D�S$0��<��r��݌�j(�$�#�����i>��} ���[f�/V�2V���J�`����Nܻ��yj`Ⱦ�Q�Έ��Q��	�ҸW�'������v*��W�\u�4U%��|��|�)7	�^�J�I����m�r�ci1n�I&qB_Wb�D��T쑊�44Rd��9 �8#EG�u��*!��mx��s��~�G�5I���R=�ޒՍj��l�^�M���l<��0'��,���X�����-#���f����s��Ş���|� �f��Tk��U����1�/�V`qd����O�Z����!?Ե�\�L�� ��b�㺊�)�0E���M�6�2�Lƈ�������S�1�� ں,�;����7H?�Ё?�6�}��e�0yJѦ+�����ZJ|,Pa���Qga�ӵ�+>1�� :hY1�%�-l����.�c,₆��e:��.B�LtnU���}�i���A�2W��m6Lс�TEO��\^��G��V��8����8#2����x�B�)���;q��G�U��^���~������?&i�W2ug�)�ϖ^F���n#��?�����'Y��~��$-ĉ��E��#�g�H���-s�H� �b�-趾�|����(�L16