XlxV64EB    fa00    2e00�p�������oZg�O���$�y������_D�ёu��[ݺ�~�'(+F�J��˶��oB���@W$`�r�S��ְč�����&�,1?%\ Y�2-G�G�ƶ�]oh�U$�$��;c�J���l������dL3��ڛ�����J��bOʻ�K
J�J���\�el�V 8Jޢ��Y4vM��1�&Q���;	cj����<d �D�SqT�s�0�㯣���!�����`�2T�LP$J���VůJ(uk1���L��LP����y��P�_�k(0�����p��y�)&.�����ޝ@����{�4�ܥ����s��r�o
��\��Pmy�+ĀU<���K<߼���	����-�P�ݢթUJ� D�Ňl�*��l��Ja�	{�Z�P�y5�s�7I\lû��8�+�m�DLA�Od���'��"�r�:^��+O�L"�����05|v�|�������eG& �����'.�ᘥf�5���_��zD�V��"m����!gw8F�f֛A�	V��@��Q����W�`���߅���@|�&N�t�q�	�M{+�*�d�W�ng��ܫC�݈�:��G�������ux1Tt`6!��*Ic�/w5ӡJ"��f��ţo巸p4��@��?q}��Y� ��^�˼c����'��)�l@��\��������F���±1��jQ��5���a$���@���IU�����C����4a*{�q�!��q��@N�yNu�w�9�N\q>XH�H=B��[׺�,��Rɻ�SBl�o�RUDW�[֫6��t-z!
v)�iqbΦ��"��H�T�N��blf^��<�DI8p���J�~�@���uAA�Q���ᑣB ��4�,�u��.vV���1���\z��z�ܖmZtoVğe܍v�	mc�۲�yO��ߧ�����'��O`��F��8��|u�Jê�r�=�� ���aZvQʚ�}��ӽ�H+F&`.# �=�ڷ���^��e�!4.V2o���Z$��S5N�e��T�@�I�K���f9��k�����(�ݒ)#��0�S�^/���׻W��K:�\^��،]�DwX����e>(|i��j�oj������Cg� W�Mэ�mJ���K���Ih�-����zBuSJ�R�-pϸe�Ԣ*��UFU�ݯM�]שV�����_ů�׺J	��v֒dΊ/��a@�k���ͭ�D+h^�L�2J.
�s;�bS��(@<
�ڣƓZΛf��!2`�ۑ��C�m��l�NiN�=�=�-�yq���i��5�g�$��	k�q{���j������$�取M�t�l��b��(��-94a�#:��U�y5��y�$ˌA��gZ���$t�8�j�WW��a� O�ϒb]KJ��� 4�J�5�oj�7T'x�r]O���lz	��L�O	�Κ[��Fw0��쏲l�~�c�03�,%3�����d�憎&�vQφ�_����ݳ��&��mZt��Ki�c��&w].�-dO����"�ɮ�Q�d�EH�K/m)�*>����m��D�����02��M�+S<���o �K�b�}�6�R�H6�麂�ŔƷE���|Y5�d�x@�E�܌Rm��r`�Nd�̂������wWr��D"+�����آ�� �0
�L�#�Z���)�M���>q:C�+/�oT�j��=¨%�RyZޘhݩ����q�Y*ڛ*�%76�Q�.TW$�����d�O����{ۀ|��7O\�tj^�f�#�ۗ��tj�;�>i�qs�����W-�f�ð����J��m���n}�_I1ۢ�QmO�=Cv��N�8��D"�Da�б��J
�mE��s�k�kpun�c���}�\he�����^�NAU�C9�%�U�������KΌ3Hs㯠��|ݧ��Z�?�s�*�bS�%Ln[h��H<�Q�y�y՝�#:�	�1�<����!��c$~=�ۧ�}�M�=�+C��L��V/	���Q�9��;��(��<ꁜ�Ċ]Z'V�`�_m�U!\4D2=:�z��o�[����^�OG�+���Sy��2�{\���L}~����������e�L���@�?1:�V��~�q91% �˂3Ĭ�I��Aq�l*�u�s\��w��ڥ��tPBz�\�~o��-!�Y��=�����;�:$�Έ���c(�ƨg�ZM*xE�����#�CK���+�L:-�޸�Ӊ�!䴗�c_,�Yql=pL��ӥ�w����I�8�����D��s��/�J4��&����g4�^zY A��τɐLx��9{������pޟ��1�D�� _./~~ͨ�f!�YaQ�ޛ^ G��������N ��wY,ӂd��� ?C<ʔ�a�JRy�u���2��Z�hWs�R2yWYS�7݇����	���[�,��tc�~�8��?׍}��v8P��&��vɆɟ���es�� �=��ˮnl'jF\v��Klb+w��nj�q4>�Cb���NX�:��2G
�띛��J�<8+l*ϳhX��S�-��_�u�O��Y������z�����5��Su�V��TmC"�H���M�d��'���0Z��H^���=\�4�b�M��X~q�旿�9���0�˹�צ;'@��i�i&l����ޑǅP��G<�̑��p�&vF6t-}�������A��p�PT��F�O:�x��� ��{Z�T�kx��.�G����|k�
��$����]��2I���j�1%ȑ�(��<x)�~Q�k2>R�&�Ⱥ��o-�u)��0 e:n�����|:��+�'�������+:��D�_L�a�#�'�ûyk��^� ��-L�i�O:6�g����)���,�"��w;{(E�f�]����d�T�Zd�L�@�V��Q�upI���:`����Z����Uxn��2�
c�q��ݟ�4���9��n�a�݁8W<�ScH�r��7�L��Wr 0��5t�_�ӑG�z��F�;V�o��u��x�oT�͠#|`�W=\���.�{� ������//�� ���������a|�o��K{!N���;�+@�؅	^�Y^���g��;S�����������>�����ĝ�mt���Y��	M�c�d���%%��Idk|���ջ�.b�/#KfX��nP��'?�a�Q\�5f�+�Ԁ[��e6Ϝ��<���(&��[�c4��Q��bo��Ep���a��3j5UĮ�%:ed�sCZ-���(�:��,P�Ԫ����E��P=ݦԝ���E����=�r��$Hr=�'O� ��6(Vh<�Ad�A+�����̾��텮H.kiua�J����ʧ�tچ���e
����ѧ6|�\�Ea�Q.+�R����$��R�7��sҤ_8�W)[���D�5��~�)�?��w�ڃ�/u�ڳ��l�e��aY�Ӡ��/�m���;��o�2)�k��Sp@�ˠ�?ӧ]���cɲݔ5�)��$&�Ӄ���2�q���E�6�p�.צ�?�_�oT�~�\���=м4��X�Ah?&��k-�oq?�wg�t?��k����ޑmM����q���[�͟Q.KsH*�{Ԑ���UPZ�(���.K�͑^X��-��Xq�_�*�%vvPyP���(AeE=#��Ym��^r�&�
K��R��m�"���8Hs�	3UW��SB����'�����Md�{�R��IU.��v���,`u%�e��e�I��k�A||���r�*\�W�(���z��:
���Y���-!�z��i��
�2[���.�H7�,�6.荢$ٓH,�y�Kx��l��԰Ze4�uT:	��&m����t]��Cu�i!�Pgد	xf���Pܞg�˰*?��Ȱ'
�(K�;%�<f/�T�dwu]J/��>�Q9�5�Y�WZ��fgM���!Ql	��>ٜ���*����K#��$��=�FD�m�4JT.EYJS��������s�Y��п��v/vW=�Ł��SC����8�>F�A f<>h��a�-pN�`eH�bxY1���:Z�a*`�' ����9����xQ���&�N�;�u!gB�'pϴ��i6@��~A%-��:�= 
��6���c$h�韭�7�1�US�S0����e�z֚�w/�P}���[6�ڜ&[�	L��"��H�q���~�.O�����8ܘ|0�v8<�ȹ��7�N>	fw�⢱3\��Bz����R�}�]0��+���&%&zzQK�zؖj�r�E��"�I�P[@����=}���\G 
�ZJ��s��ŭq�b��O�������B��>B�J|��s�����X��/�ȄN2�/���
��v�f�/@f]�r��	>�z��R=�����F�a��O����/Geߏ����E/K]���xyK_,�qK_�y���ך�jT��Rf��~٘]�&kk۾����]�Yu�S��!>�4��}�D���-���]M�3�Y�V��CZ�]<�1]��� -�qocÀ�7رԥ�B��9�X0K|Q6>�p�5zS������A��*�HU.�3j|ȶ�z�J����Y��t��ߡ�p?`�t1�P�
��A�d_�{���*l��ΩABn����S���� �N���-�@>�z�2N4|��
��;
]��\+�%�q+�u}����W��Ll>P�֮����2�\|Ic�����`�����r�(n$�!�iV��E�2�i�l���V�֥JI$��>cW���*-.���8�4Q�_� X��:=��4j#�E�)
�%�\k�|�d�c��&�� 	�F��)ۊ�i�~e�k�>�|�]�5;�h�:�z#(]�`��$o��v5ݵc��ߍ���_�v+Č�UX����!B�aC�Aq�je�Q��#)}��SW��v9+u����g����z�����*���n�е"N��.\h�E9D� �^�a���1���]N���fz�����7wE��a�"�^c�3Ad��T��9Z:''��_nZ�j�a���A�(O<hޗ��m�<rѷ�T�9�"�u����/IZA��b��`P��a6�K�1Et�)��O��@�txZޝ�c"��O�)wܺ����tE2���9���Ҷ��u�s�w(�&}'c@�p{"�!}��[�Ӝݚ��ѻ%F���§Tș�/o�IX���mu-�3A�2K���?L8���bv��V;��l�:�� �_��n�oyW�>�6-iE�L~����./x)���J/��+8���M��p�y�I.9�
�������s���&�K*0"!����mBs�0��ɘs�i"���@ybN�
�=^_ldT�h��05k[���m6Q��a.f��O�,)4����=c����!9'�<�c���<+ZN9`������3�E@���fJ>(j�@w���9��:���
4�Y�~�
��\��3�{N6/Al��r��i�y���>5�u��ګ¡$d<�ddMϟB�JE,�eع� n(+`e|�����Z��U��ʗ�}���g�e%��j�L��9��i9���'��'fXP�B3��{�^l�.sB��g����ߢ���@�I��6�-�D�1&EJ����6�p���������i}�髲�&�I�≙Ƚ��_��ݵͧb�&3aa�3K�qXd����k�k莥'C�)V�PI�;Y8Y�х���a��bA ֙!�0��^���C���_�6
V-(��f9c�s�~+YTs�xHeȶ��$�|�Be�m�2g�6,&��,,Jl��6���T���6��Tt�ACd��B���.[}@Λu��/��&?i��G��L)W�����'�3AJ�u��m����3Dh�L��c�#�jf�*�0�[�>T�IM�ɷr�<���w$�P�/ёῥ{�a%������j`v$P�	�����!��Z� �����a#����x6	)T�r�.&0B�x�ܲ
�:���"8�0�Z,ם��"=��e?���� ���6�W���#yue2�)�WI�}Uo�,�����L
{tQ���l��d�E�T��\<F8hlg�F �Y������=��~��y"���|�#t-?XK�a[�'�A���#n���%+z�'����!6���B�2G����>��o����[R��#��P�T�D}�"[���CF��Դ��<�=�F���ĭ���s�ʵ$�j*���m��}27+u���?*����7^�U��ۅQ��Q��6�	���|Ȉ��T+�{�8MH�c�EWI�ۢG{n���B�F�c��zi��|e˞'��a!Ƒ��N��5�Fl%�7��� Z�m��SZP�r#Ն����4}r�7BYu�������!�S�e�,�*�C&G�&��D�#:mXGѯ�1*h����z��ۇ��VN�4������SQ���تM��\To�1#�P�Ft����k�ҮfJHJ�v�f��6�������6���o��ڮ���4�O�9�s{��nL8�UBxռ$TQa�	��k��U�1�M�b˶VN
Ӆ�����}W;,k�kPy|ɶdd��K����9
q�.��zz�5��;l~���~;���A�5Ǩw@)��1��}�7'�R'kE�|��N
['X�2�x��k	N���2;>�z��y����[3�X��&���	Qa3(�d0�F��Ig���4� '�f��
<����� =�n�����r��O`�,+�`�u�.�-�^��001�55������;�<=�J'�\�QnD[�&j�}�>�jl"�|�F��&��ͧsa��Z��4�w����ng O�w��J4j
,Q�� 5 fv�݆���e�.���Re�j?���������@q���Wx$��$'M8'rj�	�Bs�P�����L�T4�c)J�=4��D���` x�,���k;g�r!���u� Q�AC~Bͼ����(�@�F��ZR��Ml'~��M��
6�pMxařVP�VJLߟ�˂�́�lw�q��.1��SϺ�TRJ��KC��x��5ض��?,�&p�lN�?��� �!y�dLiC�`����f����\�~��TY7ls�ͯ�!���eG����.D]�t{�{w� ,�v��p�%Z=(�|�I����k䇊Ej��ecޣ��Z-����WZ~��l�iw��*N�Z�L�c<�&���fM��=��v�����ީ����F��'���򴞨:H�MT�^:��蓭��p"�y�����'l꿪�P-9fxH�p�,[u����g:< D�p>q3�9�Ϸ.,^-�0[��T����p+�ț�9,�Z���g0Ϝ�8�Nư+i~�-s�佮)��E�����F��DE���#=��13 �3��Ki���g���z�?����nk�{����C���L���$�BS��d�f��˯G]dsޑ��=ޡr�Ͼӷ���?@��Ħ-Ȗ}x_~Ê9��.7�X67���ٔ���
�W��:F�a���t
D�YQ�/������K��Z�b�H~k�Cf�$ 6�q44�=ȩ���u|@u�,l��ι4�F�
-�9��Ǳ!�_�ߟ'��{Xۍ�2e*��ҳ�pky5������ʚс�P��W�\v�-�r`�?	lޘF���\'<�&*]�0VD -2{���k�c�R��0C�W;�QX�O�V��I�U����O�N	����)�:�n&ZQX����w�����^	�z��	��tK Ͽ�G���|T���_��4>UC�@�j
͔R�`�uK��!'J?�cm��(��]ˣ���q�W7��f+5xn0O���{��
N�/��}g�X��A�^�>�+�y�3�g4�YӬ�&'kh���4ڍQ�������^���7�$S91g|�I_C���ޞ�]Y ��)�8~��s8c�A��T�q�ed�����o���@K7�Z�$Bs֕��� jϿ�C�	�A�P�V ��^�ԫ[m'Xv�9���N|Ivf��EBk��Sj��l��g�>鍟f�E�e�x�Z�'���8wG5�c��B���EzE �h�ς��]��mU�y]R.���yN���1�7�8<�N��]� �%�j���n�HD� ��L����
I�I�ў�m[��Y;��7/�	�Y\�M�m�*;�`��)3[D����ШZ��%�Ox�<O�z�C���`2A� �;l�&a�$�l�����%cT���t	��ʡ�3��E�ϯ&Z��� �4����?";�952u���㗌���ͰǩZ��N^;�l����`��fP��j�1�7Eg�X���[_*eU�L���D�r�4�|E����Bf�ˊ�GW�H��O��G�_OLD�f��M�U5U/�R�$����b��$�n���P����B�){�$1u�.���KH��N�p8|��ͳ��@:���_yB �\xp�p�4��֋�����q��5��e�%.����)m�We�Y}�;������؎p\HӸ-���-��ahg��Lfa;[������_�'WT��m<L�<uH��1���?5�`�훺۽��J47��ؚO�+>���j�$D)w���S��V9_����b�N���p�s?Ef���]�u�ZP�7���k�h�^�7�5�8}���Q^�刘@���,
����)&��a5�a�Փ�j���ü�A�M�x�Qu!�yϰ��G�6B��9Γ���iG��V��m~��9o�UX�Ae��<��n����}<��|M
V�)&r��i�k��O;��Gv�m�Z[Y�N�[�*���(��?��L%��y�/��u=kA�&��A_��\�c5�v`� �e&�8�WIɿކC!Eac9x2��2��V,�5�� �����NEW���nzaf�)6s�*Κ���]�c����Щ���RC�|��'�N��O����ɸ����ҫ��^�B2�����6��� X��\�GyBh��}�)����aS
�
�Ƈ�s`Ý�l>G: f���<�4�;M=��|A|����11?����'q��^p����fs��A"8���Qu�,swj-�x�����R���������@<A���?oٞ��B�Q�x�*�b3IE��l�`�����0z��է��P�]��8Q�k�ؚ6SC�9
�'4fD	�%�ux�nU4z����z�;�ǧ�Lz�{=r�A��-#֐�U��e;;��3� 	4�=ʳLոWʾ�$sL}�nן쟗�vKȏ�
����"^���#�U��7����j����L�4!�e��T�ɿ�Ŝ��v�[�����$+�e�� �$A����t����`<s������L&5#���<��������N�Y�<,�ksM�&��h,��^1^UI�}�6l.�R�yZ���OE�����L�s�ȇ �qh��o��䐸�?Ԯ��������"�1_����ӹ�L����Y���0V�lC/��6��x�Zn�L�M��U���&l#VL[F��!��&��E�,�=BPu6-������۱^���CO-lg�����L�^�,e�ڎ['�V�E�!����J>l}�6�3��nr~��}	�{	�c--edV�;0(�G�����$f#!�Hϲ��l텃�Ld�����w��2vIXz��` Ty�����^8�o���g���������pC�=>�n�&�;�9t��N4
��Er���+@i��'�~��Z�z���S��
���b�? �):f'���$ [�F���	�'�<a9��I��<4��k�LJ�ZvFi{M���RT)���SD�fdXɭ��}R�s�ӶZ-�E\�9}����z��NM��i^|�$B��>��'���|�>�M����*��}0 ��%e��9�b�`�I�->�Xa�����c C,�I�>�2z�Xa���l��"�O�=��+�T�y��9���1I��5,�6X���t��{�����%A��;(P����*4�~
)Pv�I=cG�J�Q Q��_���{ld���܂���Q�Z�5<��#�Fv �CW��}1�w���c��s�9r����	���є�9D̅�6����oh���T�Ǧ�$!�{���^@�#�ct5ޗ��NF���Bt���p���{��_%��B�m5�6�TI�a{���p�\h�ݥ8�Q�p̴.v ��Z�&pa��S���	��,m�l�f;y>:�8|��@��B��f�+�{���@��揶�E:��6e�]�gC��RPS�}y�g,4Kݏ;��6
�"u�Cb���t���G.φ����34W�����嵌�=� feR�>w��s���\hA0������N���"�㏦�oG��=�	�ձ�R6��h��"!Je �e�77�~���uԩz�BK/���zB�.95m�vL���M���p����Kd&��'��7��I���R8%FJ�zN�nۓ�?]���HE�C��1�0������#~��h��q�	
U.�?���{�?i��0E�DK��Ho��@��D=M�Oe��?�'���E�L�u�"t=�RӁ��@����u1*ƈ�7��/����ؚ4bD���]��9�dd���6�o�`p	���a��}�E� b
|o��� �;w����hg����;(�BCa�g��Z�{?U:����S��y��N��L��iV���f���iY��:��d��hJԪ��Xj��0�W�<��do��)OFT��d�v���>�?	�;2�r�9�7�zĂ���W�4���1�0R�6M%��br�Q��g�-x���ٻ�/B���Y��Yu]�����|�2�*��2j�2Gax �''y(�
��6+�	�6yvT>�Ҥvk�LE�	��+{q�K��mOh6�Z���'�6JҀ�A����e4(���"6��)��ZnHv~�5�\͔�S'u����"�Rm�`�"��U5��A��� ���d�]�qn +���d�B�<����_oBC���d�fMmwY���x����#�i�6@��¨�U��7��E���n��!�Jn����Q��@#~�K�7,�4��+�y�(O:����]ڵ��$¯��f���<����;���y������(���l@Y�ח��^� ��߽�*w�~nqʭ��'�������0m�����yٍ���+r3P;�����{X@�Q'��R!.���6֒U�es�Y��d��,�sՇ��x�C5���X�9f&
4�9����6� :s.Bo�ew,`.��7-����-ks��jY�����YH|�Ȥx�&uV]�$�5El����=�}}��Y=l�`��3����\���~U�Q�:��ҳ�F�n�E,x�3m��ْ_����Oe_o����a	��@����u����Œ�8	�=2�D���KS�i��թ1f�G�~�,��u_T�pZ �fb��MG���J�Er�9W��:��	��������
K��BEm�*���;1�|`�h����u�g�q��dB j�!��	��Hؿ+�9;��P��y�b���������Yo���J�{�O�3�XlxV64EB    b353    1b50w�\�3�i�섴�r(?��rƹN��z����{ӘH��㵖�7�����@��x���:g�5͑�Ajz�YC��"NY�f6�O~4YE�����.����D�f��Hf\JC�yJ۾�����9�4�_nh��,�9Wt�E��1��re���8j��q����Dc�&U�6�=��ҫ��x}_����=mۡ�����ʧ ��R���C�}B w�$7U0���Rʩ J��~��뢞�`x��oo�ѽrF��Zz���������e�",��i�F����wb�:�g_�s_��l׉�D+q��݉�Yv��t_�������)�z�I��ʒ_�����8r]���~Da�|�����	șݝf��1_M�H�!�&�w���}>W��Պ6��=D�P�ēPr"%��&x.��`�!�C����"2�a�]m���vV3�TPq��	:�bsv�q���?�e�p&Wha.��P������Ѩ� �����������$�Z��rS������g:�#,�(m/j:Z��!E{��V�u�voPQ+�"��FF,~a�i��q���������r���P-��չ�^��8�!<v"�"K�X�kQ�2Y'Zҳ���!�I��ƫ	h��G�1���j���|�D���NQ�I�����GN����l ��5SI�%��{������ͼp73D����n����_���ڙ ��J  _@�ۯ����B�;��p'��nh6x4����# ���ޜq�U?��݉�X�y�F���r=>�i�g��(U���O�Af�Wgv���c�ޞ�X��\��ɋ�K���a������P\V�כ�s*d��<︎�����}�_ul@�Q�����۴1"<��I��^�>��������l�Tn|���tV�`l���x�W�@�?�c��,2P��G_v%ǯЎ�#�E^�|R��M��J�3׀[�����;)�?�)�)���|�g�S
��U<�e#y8�"�1,��Y��2�@��"�7��o���\�m����������}�.�Q��e0g6Z�+���,9]�?�M\�� /�Bx5�$�5|�N~�On*�(ܵo�?���y����#It8�{K�|���A���wXZ-����Α�|�ޜO��C~�`�;6=���1�2~rSmń?X�[��p.>]1���RA�J�,��T���٩o�n���vO���)����&[E���l?��hU�!AŶ��]�N�+k�;6`�lN�zB4G�a��:eQ1���R6�,�H�������3��e�	r1��T��g8�X���p�V���?LMp�C�j=&h!_]]mƭYj|�佞�����5��߼]�2yj�`����W��n)A{���$�x�����o�^!h���*S3�O��;
u=6�Hh��6�Uߟ�$Tv��uNv!��)����ܷBtl�M�X���g���=�?�2�~ol�%}��C�Pv8�� ������dd�Cp��uo���G>ǈ��ju.VJW�a[��5b%ђ��{<m�C���O�?,T�@y�ʇc���o����{F�wo|�����^�}����w��~3��_�}�8����@i�X�V��&��UXZ}[������@�:`�`9�]�8�.&5=�-�U����z/GPO9W�t�f�Շ�4]����<J;��`g��ɥ�8a=�
'H������|dSD,�$���i��s_��D#5�<X�N�n�*�r�/�圠u:����"��B�_cS�w1X�7��S#)_M�YF�o��A���3�_��i����Jwp[�ȬϠ���S�j�*{�u���%�������o��-IQ�^�p�;>瀄�^YF�rC>(�8(�fZ��i�Ѓz5�I���%��j��Y�:e�_�mI�+%EE��"L��X����y�W��N���S����S���P
eb�E�R�Q��������)�!�_;n��/�z^�WbS���_�ӁG���y���r:7v���R�92�	�66�Că&��]�d�8RP�H�?F�Bc�������c��Rvj��(�z'�Cߥ/�
s�o{w_����>h��(������j�S����fN�����~�X P�VY�"/��`]h3a�u��ɴ���5����k����\�_��oJ|QV�w�ܧ�����i�!�b7�����Rl˷����`u<���>K��X�Ee7�<�ev�]���8]�}U��m��SLCQ�Z_��Uu�F%�U%ׂ>>'�����.}��^|d��ޠm���BTR ׯ**6��Њ~L��,���bR_�)�6�F0N(�N�ie�ܿ�-��0���WHm��6�`�y�|�7����(v����N.m�42%͍��^,����!L�.��OZ�|�h��a)���Ϣ� -0��?��ͧ�5H�|�_��Nv">tsu��H�;i�:�ΖI2̠� [�YS-c9��ܺ���P�3l`i�5,$DV�S�4���P=掋���Z����q\~|_i4�߯��3�|�4Q�G��ܩHs���ػm�y1�l��#'P܋Z'�)�W��{�%��������(���$�M}E�����wG��>��d����&���i\�KH�μ9b##�E�7j�������T�ΦP�����
�EDt�Ft��{�¡6�K�TRu���E����6���RPm�3J8X�N?$��X��6 S��'����TMn����b0ޛ�
a�|zn��n����&s��yH�v�+S��4�����Jl�0��ө���[�<ќt-�!Y��*���N���S�0_�36�����) �Ov��r�I���HY;��ގw�]46��[�=��Vm�V�;i���'�R��'��j�d��
΄��Zc�o��u���r�`�)�ӭc	p�����|��*�#%�2�m����I�œ�+ϓ#u��td�\q�vB7b�9
�[���2��Q�:��u2jژQjF#P �H˶��57-s�[���Z}F>m�J���s�����ܹ�\Ş�-	�]T@�?�� v��| 9ɱ\����-��>���;�4�hg�l��� vS(���)�� �C'�e�UZւ<�����>؎F�c��E�G��j���\4��H }�HU5c��M/x|ڤ0F�"�<�^�h����!����������ȅB3rm�7b
�K|Æ�C�fyG"��hm1qҊ�"\ ����2��� ܻ���ۙ�6{�9���}Sk��M��l����n�q#�R�� ��QXa�z~���:�A[�}��wq&���s{N����X�Th���"��]���*S���%��)�:1�U�	�,4�"�b���[b��9��e�,�F`:Y��h�͹ ���༚�����h�e��6I"KhI��Ñ�Tw�H�Lcn�� ����E�?d u���O��R�qS{�iN����-�=��b�Q�{W����9�X/lr8��*�G����?��?�X��L�p�8���bӜ3��B75KJ�E��]8b��sV0���X���㫗=g�WY;j�y���y��Y�5I����'Q�JX�O�T���'_��v��Z�X��i	�,3��ֆ5fF�4����~7j�|y�mP��)ž68�͡8'�0J�ןQ5:�?:R�Wg��D��`�n7���1)fY^�x���P��K8>�����HS\����o�n���w�n{�wm�S��h(_)����	b/�ѣ�D�����6���δ��@�� r�e!�4��?h[���S�k����|Q����Y^���&Vm�F�S��ylhmBߺ�
���@��$����hQ�ѲbYdtJ��4G���`1�?z��t�fy�w��Et`�R��~P�R�|F�jg��y�r�?��\�8�:���p��͈��=aӑ&>�<t%�$��� ��S":Ґ�44���a%�6���ذ����� �V��
�
y3R�3�^��U��F���v��n�.��u�'B��J+=��'64��S��r&;!��o��W��G��|�Dc�4�7k�Dftm>���8̴v�2dGs�_�H)^i�¡��0���єKQ;R���=Ҽ��� �=�����L:�d���W_uy��oP��4%>	����c����U�~���r�uηo\s&F��Fc$E�;��˶�I	o�����on��(In>͂�����T�i6�۔�4�E� �'� RxN��%�L�֠.;i�=��wB36���nl������������N�"F�i�'�!�b�qe#��hX�Ⱥ�yW��V�a�<:���1ՓC�&�d�Ig�7�=�����4���a2���tD5��B�ed��m:hm$�+
�$��/X��ј?��Yy��49���x�Y�I��o��̉b8����d,1at��=�h	Jh�f��S|e�+�����Ok�z�WP�.F�ҵq�Y�$�5���ʩ�ڽ�ǆ���P+�Y��g�UP���нpj=�#�pt��&�&����m�wn��
L9,
�"ʀԓ��*?���] �|�ܿRm�d�f�yo|�j��{�`>�tu��Ur�/��l��}��w��;h8�X6d�;5��A'��������f�ߤ���!��)�o&��͂���J�8��J[X?M!���aI�lHc5Z�0�\�#}�JVWT7 �"TW�@k�"�9A`Q~�lvB'b������
����{�`�����^i�_�Ԟ|�k����"eo�����]	Pt��8U}M�����X��:�ҷ�N���z3ΜS����Tl�:`��Ⱥ�]�泄�6���'('�ũ��B�h;�Bʧ�^sՕ��_���VRr9&(5x��#q �����1��^Gf���d���ܨ�:C�d���]��b�&�^���"<z��~�x�*mb�!��I��?�����m��B���*�0�iV����>�5��R�W�ĺ{dG�0���%v�����DA-7��j�Q2�T�V9�v����m3p�ݷ$5�Bz�6$�'�sMD[������?^��QDW]��9��L�嬏���l��09K�+�.���Y���}��a�GY���֬+`^����SA��Z�[	���.���S���Wp۴7�����2ߚ�s󖑄)bLiO�/�&e��!�pe޸]�yp�EJ�A=Ib��x�C{�7���vҴ��X& ��GF�tuV����*2�䯪�Wd�hz�#�����_~Qn\��XH�`V��>��(=У+��OܪR������������ǭ���M�3Z��3o��EQ�e�l�+��<e�
R�)T��a<Z%��]�\�j�CC>�iw��};��=M�f5J���v��)O!�i�CA���+�ޙ>�����{�R�Ә6�ٟ�qئ�������Qpls���L���|	�agή��(�N���^���lD�򚌲mg��M��\�Y�Lc�O\�c��Հ��� HoÍdf��$�9Ph��jѱ�g��k�TſPBQ�s���"�2z[�7�6���=#o0��d�_���=����P$j�?{>�'U#N��[�ݱ}KV���un�Z��6�Ĵ#����r��F,?�7[��H�7ds6l-�����x8�8����G�?R�ƒ'U�<PD�ȭ�2��R�l���N�_QL�`�Nk��p�m�{R��a��&m�0f�0�*_��i�S��7%C�0r�t�#y�~��_�g�M�����l,a2�=r�������5��>83���.����$���<���g�/��+��+��.�"������(h��|h	�m9�f�h��8�$��j����y~,��)D��W��r����rl���o�d��u�߻����Q��&k�q�p7e��Eh�`(�-��L�q��ű��M�XxpZBz_�[Զ<Ap��$�S� ���_�p)>D���>;%�sS:K�׎�SI�e_+o�ů�Y�Q�ȡ�8�f�ƨ������$�Ń�;�__ګ��ay���WG�w�sV���$�^ �V�{3��0.�0� *����!nr��)�#׳J��c	���V���`�?�A� h�<��P�z�ۏd���v�V��Q�G�����.�|k�&���g&'6�5ch�Ϲ%)�(�Pc�v$�D>�Z#I��������eI0.��S�-�aYD̙+��=Z�G-��M�t��$��~"$�D���^ �A!Cwv%�{�(f����׶^���b���V&�+�O�
�m/��}�)ᔯ��\1Z�����a5ȳ\ݥ��H�k���9��걦x��q8��,h�Q��d*|�螛����٥7�ڤ�=���n{�o�d2&e��T�T�6���pd_�y��ԁb��L���ؐ�'H7�:i���'L �eMҩ��=p����/@�I��`.�*K�(�^ی�N�}�I���zE1���Ĥ$޸�A��Mq ����8Z�yBX�-��`Q-!]�/u�5�o��A�E՜{����x|_# [���F˸ ��Sd-1�y?]y��d40��9�����|dg���EaL/Phf�~ɓI�Y_�����v}��w[}{Ws����鏤f]��%3�}W�!�)chCa����7�Sw����Ce�H�\j���Y�B�\�i��L~+d�M?Z�� ����g�"��x��m�����=ema=���m�`�"���p�3����C��d��T3��8��Q\��,E1�}���v�S�2�7�1��B������E��Nö��&A�ksw�C�X�0��J��d0D���t]�D�0Ј�[�"�P6�:d9t?�M=2� }�TrM��0����Fb���#���2��>&