XlxV64EB    17e7     9b0��b�O�� ��z��{H���Qz�M}t�ǩL�L8(h�.�c��8o���{%t��Dթ��ּGw]� �ّZ�ʱ9��#�T��u�ݔ�컖(�#���3�Cq��Yx2�emj�8:�������y.D���7�4�9N��7HJ�>��tZ$���c�S��Hp`��"N�d�=�t>�'���%��&���t���i:���DA�J}����ZJRӘ��{��	[���PӨ+4m��n�7RK��z��l{��u[�]�oKXF�^���I�-�1�|J����Q֛��J��LU�ʣO�4��l/=o�32��G�]mE5+bd�(MB�C�Jq�41�C�a��,�=P�I�,*>�J9�#�4�ih�����@��;��58S"�ulN�HI���l�ɒ��wBq�0*����oz@ؑ�b�SUa�5�{�)L�`����NG�X,x��	�m�r,�9<u� Q�W]�}�D���_��\j5�1��X=�������IKc�/�8����F=,
HƟ=������`�~����d�'@#&�O� d�(����)Z.��ὣ� �G���g��㖶�>�
S��F��p�7��R�����7��Y�>�V�,��I��r�q�/��Q�)����O��%no�9���.ማ5R͙q-G�h�+Ӳ*��d���zi�>�Cr��)g�~����Z�O�0ǁlK��.������u\�����ٔ@76�gc�;��é:Z�r��@I9�*���@���	UM��k���9V&d�%���p%P6�l�#<	e�$�B���s�W�C�-{K	�>#���&=m��zb��m���s;0�:���0c+��p�52�O^��F�۸�X@�$i�I�9A�=w�ꈧA�dq8]��'�b�c�5ii6o T��xO	X��R��6��+Mlt��a�8Pm�B�����!�ϯ����>{��L����y������|�j�,��{��=���K���#�*-�}#��J���R�P�kz6`�>�"S�+�yLjJ�����n���L��D�8����#���#mdG]UC��ͳ�7���A�ağ8�,�.��Eߛ��|���
�[h4�`����x�t���=
U	��-##zj�v��@�d�Ro�f��d���[/z����Y��@~d~}����r}���.��O�ى��TN'��`���2�0L�+n����H��7"0|��N ���j���R�F����;�4��Rky)�feY���z�5t���-�&��X���{�S�G@P�����Xܡ�d>ǟ��m�;�V�rlå�&G:�O����g��d��k�cm����_�?`��v��б�pW�w[��
�&KC5M&}Ad�[����k:�>����)-��"���o�����|p���"����E�$��[��8����ݖ�p��0|j1�GKf�")��5KZ�S6'��eK��}��z���ͺ���+�$�گټ���B4Uܪn~ fK
n�e�rh�������Z;=N��tJ�^�>�g��;�Ö���Ah���U���5ք@���ZWo��D��e��ʣjT,�kq�n��/Z�_[|SZ�=��
\3P��#�Ƹ��,�ѝ���s'���۳���Q��LZ��%��٨��|cق��s_X��Y�2>�wt@��i����O<�Z�h���(I6��^�����>2��a�MI�R{w0�N~�p��>��6H�%eާ��6�Qo���Kc���ݽ�\�C��A�������)l��{��S]ukP -���PI����9�n���k=LgDt�Qٮ�+��l�A�*$ԩ�=����o���2%T�a"<i�R��q(� Z1�d��͊kX�m�N�h�=��~���x,���}�6���=�_ZM���O�m�^���p�1E��%�5�*��u��%S%�*�A�r���Lx8���BK��_F�b���P�+�gt
X'�A��X�K@�*�(Yz���ԮD�A�����O֋�[��a� �b^�dD���v���ۯ<G��d�U`:�JX@��R�,��h���S���I
Q��5څ�\R��|�X�_D�1;n�t�\�nN�5��}v�t�����3��_�2@����5 a>@s���#�Up���b7Õu�2_t������(�'�Rr�Nn�?��DI[]���̚>lT����<G$�]��=zm6�䧁nbFL8��Z�з�� x������8`<�����>���&����E:��a���':�|7l���<x5ƨ����>� ���D�e�ɻ`�u����97p�V��S�;h�~���)���=����o8;����Ӣn��ɤ�]`��\f����������O�1�_Z4|����0e��Yw�%^^D2[ZLrf""j��ŲG��