XlxV64EB    56da    1340�"]z:)iv��B�YQ[��zRV���=qk�c0jÆs�D��������fJŲ(Oja��k�0��t�F��5��5����6����ĉeJ*J8�G��s���M�H�A�,�����#�+Zf��}�`&���ֱ'i�e�g¦#�w�Ѱ#�1��>_i�]4�����&�b���h��4<���4�i��g-zꁦi$K)�E�9�����D�P<\��YY�/>*{��I �Mv�IU���ÿ�*���U�u�eԨH����L��?�i�6�4��T�hU�Y$��BM���B�a�)��H"}n�41�UlW�kOcxhɮ$ԫ2Qnj��z�c��H���	h�^ɟ��5�� о��W��h��;�&�5���ᨣ�?��=4N�K�dp�_�f.�d��<s�/�$Ť��Ѳ.L��v�#��B)^����$�1���]����(8PCA��Y�U�s�w(�x�rok3�4�G�|����<V*`��_�I׀׆I��矯����a>F�4�k��|�� y/ɺb��@K���(��9trLU��ե���f�%��
kJ@���q��9�T�����K��0v�,�;x�smA�{�:P�~�.��{�V��j6��ښO*J҈�*��(�+JL�����&o)��51+��ߌ%87��8����x#��2���k6�.���y�$�n�!l�B��W�&��k�o���=�,�a�9�D �yoP�A����vAA'�
�>8t���H�}��^k+�#��̙��%�jb�����Ȟ��2�XO��/����F�f�tV�/?��T��1Y7�����&�>|�%��ٮ��E ���e��9U$��[>c�N��F�P��>�th��^�T�6��C)����:"�c)\z��(d�8��@V���Bu���:�
�kmR��z�|���%��_����|�G+����\�7:��;�*G-6~��=x�y�@�3�(��w��|��q}B�;��æ�w���&җ$	y=�_���������d���q�V#�"�N�i?��m�y71+���/���IX�&l��W�&�;u�U���ƃHLV�V�9�4�/��L^v��7h��¼ŉ���p'�y�T�wZ�Ɗ��r�; ���{�@<��Yc�q�y�ŭ� �'f��4[��dN(iᝬ�&��J���� +�\�8�L���C� ��ڟ�.����~�T�&M��>�ܩ")=k"v�3��yh�q�Yy��	!�V<�M �w;<J>_�"&\^а�!I�E�]b�����QL�q �B�7��t���5�<�i�У�)={�]Nخ�������N����6��zG��������K�Y&�4ǉ�P�jy@���xp7���b�ӓ
�N)\���W�n6�|}&)g�uE��^{)�-9�I9Y[�|�wDWaP732�ߔ�4Z��F����J]�C�	Q0�u%H[ǖT���R4Z��I{^�ap&#�1½�/9�;N�ni(�OI��~���v�܍8�D��h��&:k�!��'�g����Y{�^��p?uE��?_Z�u��s>�	�_�$^�ѐs�,����H4�O��g�M�t���V��)�����3{��XX���s6���n�D���P�1�?9M� ��^��>���7ߞmzk�up{���ҝ˭�eg����G΍PОƷR�j�T���BЀ�*�Y]�hk8�*=�P-� �ń�(�;�H��k_��^1�&-w�c����+L�B�B�rOfIE	�P&���c0r7�~��X�U��k����3�P��O�C����r�sm�v�FCL��K)N_�1�j�chH����`���n�i�\�D~y���T�3o��e��R
�R1}a'�\u���G?�U��Zҝ}�J!U7������ւ�� �<�B �|I�O(��i���,h��r�����nb��CR�4��K1�E������4��D<��؃̥�:�b�$O���@*6n�$��o�1S��W����l;�+��oM�*�&�	��#�N(���^���t��5�����E{�v�W���OT-�BJ�+:��L�_�Ӕ|�o�Tl�bfn��9����5:�R��R�1��Δ�j�/;35ѦB��NC�fY!�7E�b�_�Ûrg-�������xY�`�T,H�?�7�:��aVa_�#+C�W��=~�@��:E��d�5~ʇ��|�����@��k����B@0���ú����)DU��rN��H���]TG�-��aDiwn�Q!���bc=���.l |e��Ɔ�֋tHW�6�1����gL&�N�$2��,QP7����XP�8�w�g��/�*#���t?��/4���m�a5�^�  (wP���nJ-��ˌ�bP�<4��i߫𳯮��b~�o례MNm�d����	��(:�c�g^zR���}�X�uyB�_[d�8���m���э6*K��|��ڴ��X�d�g�VGJp��  �b�hun��"���fZ���:U2L�H�����b�8��$�g�3��\o$3�{�ɛ����A'<�T� �O���3s�pK��/))�sU�x��GnA�,��w���~� >CX��݄��t�����0�q}<&#B��>=�Ӣ��n$c%��ᫎ��bef-3�
D|�N�X1������&e�����+�����j�l�>�xaД�콴/N=$8ܻ�}SG}�MdΑ���?�E4'v��:q���A�A;$�v��QRl��zAM��8�Ҍ�*�c�,�L����`4���O��x���Gwp,�s`�5���VV����i��F)~�D`�μ����M��hV�}UK46C�k1�t
|
� ���ej�O6v���~!���a��)MM?�~���\�B�2��!�z*��Gv�+�.p(��(��q���q�����O1�W�IN���ͭ:,�) y�>ka��nz*��[^����X��F���lQ���{1��$���R�(���FL
[S�H��泸���I�Y��&�x��a�I����5ETR��~����Wi����~��0���)�HLi�x�_�ݨK�Ht�Wie=��K��ܘ5B�հ�/aPz/�8Ap�xj�S��S3���e|S�,�%^�(�"��������{��SÆ���/��O��'1��CA�}	�2�qѱ��l9���;����D�a\	7pA���ӄpA��*���"7S�_\o2��M��k��6q�nH�����>�Ӝ`eL�K������b��(1���i�u��ZϺu���/���gы�	8�	_�OrS�iB�I�2Px>�E����4忼�&��u���\m�9�	S3�h�uz9���`�֛�|9���Sb��|�����g��`�p����_���'�ߔ�;*aЦ�+L�=��-@Xdj`��{t�@D��͒��"��B>;e�C*@���ҹ�
[j�k�E�Z�`�c��v�S@l<�����%���#�S�.���:=�D۷�C'���H��)F`�}�	MZ5U�2F�W���ɰ��{��0��{��˓I��t9ڞ-Ų09!
[N1�3h��z�M#���iӜt�Wȵ�6]���@ C�W��0 �����o��:�T�S(]sN�1/��5�xm���Zɂ�A[�VɃ�̫���s���������>J4��|R��2�C�#t�O!r6_U6�'����˴��\33|��t�췺�o��̪/H�������ڔ:��W��%�j�+��ܭO��Je��V.�ak�&X��ʹ�.&>O���̚�n�ɜ-E��gP�r�:�X59g05
�Kj������Q��حn�u].��3�E���CbS<�'͝��2n�	�>�E��ax���ɹ�8,��'!���H�o�i��#�[26��(l�('�|��Wm�u��a7�T��|�U��_w$I�8_�^d�ˢK�/��ŴF���
I�#S�(? ��O�i���(�ˬB[�+����g��w2c,Ӹ� �aS�Y����Z7|i�=�����"���%�^�²5h1��9��\��w��O���V)�L�f +Z�$)��M1���O-��f�RH&��Q,�|��nWk��l宪*�f|�V���M��͡�4gt�m��~)����{�����vp?���t��@YKX�z�t�.9�)4��F�^���?����"�$`HtN��-g���=B���?k�'r��-�� 1�d�ViQ�h����$���M�K�β4�����K��)aрńw�W��
U������/�%#B�Qڈ�)�&r��)�����@��ͅ�}'WM`���Ȅ�P,wr64�F �gP����/$�'�J؂�$���6xX�����\Pha��I����qL�c/a6V�d��fݩ�1�F��v|'Q��KA��"`(�0�э��E�f�&yԅ7�=����C��[���C��hO~áM�Zq+R��1HG*��HX
(v󃄭o*����]ޏ
�>W�w�K9	.j	�t�A^O)�)1u7��<�,�}p��Z����,�/���������P����qK"��&?��^�.��U�]-��%�y|n�؄�`g��2��v�	��}��E��},���c�^���!�X�td��p�,�ܛ�R��V`��It����v�fR�]u�q���`�U��_�ַ�C� !H�h��}��fe�-�bJz����:D�O8��������2�'��#]zs^zS�֔5%�PA^�R��_��A�xd�&�"3 A���e�avI���P�SHV����u�G�mT���e�vo�EZ?���^D