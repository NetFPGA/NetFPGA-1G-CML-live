XlxV64EB    fa00    1eb0)��d�_b�δO��/o ��~��U:���~�Ø��=lM�K	��58�(�GR:��d4[�_�Z��ra�L�J��9�Ȉ�!_U, Qn�u����8���УBEw{*�7�pt�� -�Ȅ��x��xy_��<h�x��#ݍ}���O0ēK����F��i{�`�=O9�/���Pu�s�-��^�� p+N�_���� �1����՗0��_��S;��-qi�8'ɛ���uV
�QAP�΂8�	�ݔңj���0�߮�5$|������=�����0:�vE�F9w�tf9���>~���g7��n2�釩����l�)Bȳ��C]�V�d�vs~3���Z�S�����?���b=3-q�;.�P��4�ƻxw�NT� ��M,!w>���D��ݮ��K:�;),y�N�M�B ��_������h�47��X7&���U�bT������ʽ��n"9���S�_)7���	w@�q�e�CCqF뽘��v��Gat��?H'
�o�-?����X�Ԉ���kmV�z>b77K��"�1`vｰ����6)�m��b��AHʥ1��������܅N���&��Q�ZlZC H&/�>6�1�Ę��X�okS-L<r��,��ݫ��BN��)Ew+@��3 ��d}�F5�����pyU[p���;�h{V�0�Ly����5_�J�m~�����D�󿾀3���8����vG+$I�!�Q;P!!ɂ��װ�zu�+:��/PGPD�>�����J	C�/9�Z�1�n����m���q�Kr�n~Dl�4���E��� &�Hв�Yy)a��~.:ĭv:�UL�}�����p��3A��x�~}��\����0E�9�<��G}P�rgSI��'գ��q�.���o��v�n�d�Q�����Q �"�����A�7���2*�\j�h���,�N�o� �������[��'����`X�GA'O��!�ѿ��	g��'�}$GCvA?�q)�c���y�2h��udԚBϙ�|�RM�Gƒ��Rs�]׭d���N��pڞ�M�ndq�qB�lp8�85������`��~s�ի�[*������,"�����A�+Oh8��Z� ���n��7o�0��+��4h����5d��<e�Q[���e8�3_�,Ƴʎ��%��c4�v�K�4X>����"g�Iz����.P0�O�?����M9��c��}7MNx�ی@�E<��FZ�͟�����2HҔ�pĔ�`C�	g�z�y(l�b����4�Zq�i0s6�h��	�rm��|��nx���-1��$��߀�}"��ʧ��L�q�C%|V�5��85;�7����g���/��D���,��<��	j����m�װD��O�'R_5�K��,�)m�G6Ɏ�!K�#��#��*�Yj{�~l/�(<Vچ*���x�Hp{����?`�v��hIն��O(�����#�_��d�QWbq����� ���I�s��"�@=%��P�^,L̤���!&}`�D�s���=���o�~�ܭ�WA�ؾc_&<wE������;i�.��o}�t�2�����H�&��\���#���w��b�V���ѥ� � ����͖1����梓-�8�$#	[�lgF���hv��!����Ο	��B�k���p�[0��?Y�Vc��j�R����Ϋ��#��B��<U:���s��D?�숺sI֠!��DeC����{�əM�EgO�#�k�'�b]�@+B���PX8�h���gG��`���Q�K8���O�P�"�����zp5� ���`�#��lm����9�C�W����]��Yro�C�5)(>	�f6�J����R�|ܽQ��Y�Gc@1�[Z� 
�ǘZ@�hT�P�K��H��a(*��k֛kv��l�qː���5�ƨ}�""`�Ć�}�����|�t�x�M��j�q���w����c �
��)ʣ/�����=��J6&�4k���<����{�'.�5��:�-��<��NѲ�����?�6Ny���NXf>��J�>b$^r��p?�N/m�4:D0.>i�l$���h^�?�`�e�2�ڳ+�0�����U����{2���`�U7" s�0�>��i�� jp�dǑK�"�� ���,�˅JA��D���;�hi�-Ȯ���4�T�7� �f��cCX��<�{'x�br��ݮ�U�V^��xr�4���YJZ��W<:�Kv��_�2	g�k����}S;�e���.�2��EǮS��mT�ش��_O�L��6 �~S�8���i�(ښ��:�!M��Y�_N~�W�|9(n~z=Zf��Pg��GtI�� ����[x3���
����ծ��=(�Nf�:�i bjPܵ�j�1|���gf�:{���z}��C����X�����ض`0�{�7�HF�G/,�*������{�*/D��M�nG_����*�S�n�ѱ�̋�s g�x��.�'!��)�$YmoM��e���o�>B�O�ωl�<���)
bx�7H�0�V	|��S+���>��z������0n��h���yM�̣o;��{%�流�w����&j�]��[~Q�W���Vb,�m��\ŇI��-�ƛ�&���ϭ�H�z��р��}aU���V�Hɉ�x�i]�h�k������b���������f���¼C|����&@.K.,u����bE�l�އ���3��j�<JG9	E��<s嵄�B��o��*�;�Y��ͯ�tŪ��K��;%�����aZZ��vnӁYt��>e��ob-X�����g�#o*��"�@C�!�6miW���*ͫ��q?�^RX J���g�X��E��8Ԇ�#�ʂ��u���"&x�Vֆ�����j���.v8Z9Ӽh���t�(7�N�Pd�a�c��i@ �F�=��Dms2����p;	q9y��2$.a6�B��#���Ţ��H����Gƶ�B&�c���֤ei�üǵy�<T���i
uTm�&hqjj⦋	y��nhf��Ù��e�*�̌�yl�X���9oP��e�_P�Pn!>��L�����I�C�~qFy#�M��$/��[�K��þ��l�s�)����m��4��LaZ˙vהE����,ᤸ%��Ik���� }�o�|��fP���yuT�Ѳ�~������X��)ߚvp�[#b�44�+�N6���}��<�9�RW\κM��x�^g4�QC[�TT�*�D�W��>�3-��n��E�6���v�r��L������V�%;+�\aL� r7�kC4��� kC�<X�YJ���[3�;}���D-�a�Ǖ�l��#іRw��U�J�n�s��R���}T�{T�g�N���,Q�w�
��f�%W�q\���	nD�HR�T�tU���{o�;R��	�-�ά?䉇�!q�G�K�mM�~N4�'�Y�h 5E�^ٸ0�4\�|iPm�\@�|�R�i�d������� U6a��P�x�wf�ɖnLiH`4{~��W���m!(:�W��aێ'��d�[��:QT1�/�:�t�M��zB��]�p�E�H=H�Q6X
�+�.p+Խ)2 ����컧)�ת-�^�z*�,���j��9-�G�v̜�(#l�ʒ���&���6�x�{{(����$�,�0qv����b�q+R�VB(~+8B�_VR��W�j�M(��Jj�����ʪ���|�E���ŋ@�]�UB5�:�KV.<�fG9g��"��T�EԵO3k�p#���\�a����$m�I{�����1��n�&�Z���=n�Ϋ�{S��ϊ�E��� d`��IUڛ|���t�x��x�kU^V����k�� f�Öf��u:.04��q9P�J~�BL?4��խ����+K�?i.��t�RƤx*4�|���ׂ����,\�_f�>�m��Me5�d�Jq ���K�#<��&����+��N����/���[~c�d;�T����#@���{0��/tRaoȤ��w�`��ޙG0�q�����9���e��܅\�V����Ė��X�ˁp�Y>�̀�V��ɠԌ��Hj �7uw�r`đY��Rꪤ9�;R�Co?�ҭ��g�Qk���(X��r�Ζ�^V(H9�0N�Ir��(�v��7��j�(d�o��>�M�����:X�t�xv����k�?��P/��֦z�講G:O�MMX=�R�3�@�pSڣS��\�fz碌�xIQ�T��P�'|�BG��~���b��0q�:]���?����I�a��/J>W[�s�~!�O�L8�����Ǿ�{�*mŁ.��45c.FT�&�q-|u��dT�sA���� @�Tg2�KK%�O��&.���`��g�B�P̺=x�������x1��}�1��{��	l�^O��7��9]0��w'J"5*�9 �Ư�X����}����}
	H@�������į��S>U�=���^���\�،�G�Jh��2�
&�,N`ǌ�l�L�dp�[��t�i�������hE���X��f���?��7��+�]OL��av3��?��n��z��P繋	�o�D§K�zT �����C��u�\��c������|�d%2�?�y>�����Bb
� ���G=��bu���'�׏�^bj�\�+�aC2{��?Z�i�Yߒ���0�4���Y���5Q�!�ɷU��w_�1���4�M����9�."�)Y��(��M��qm	���Ƈx���Z�Q!�o�����E�7�Fd�J��C�N�{1<����a*1ī�mŬ_䔉챼3�8չ�`��v�ǸN��H��n6�=���1�v@V�-�D_�05�#��Ŕd� ���B���r��BZ�9�ʝ�j�D��X�8����]˳[_��0-����Q�"�X��4��c��Y�|�=~�V�l��Bw�wUV���^om�a�TƉ�3��j�b�65ej1�&�RK���7������+�U{�V�x�M �'��"�d��N�/���X����,VM�ɠhC.Հ��ܻ��[Q��6�h� �'6X�OF�3&��r{viX��N6���L��E
�!�|)���W<��k�'o"Y*���wIU�r���L������2�4� K���}b��"U��E�;�"����۷��L�|6��i�Ôy���El�7i�i��-�J��dΈv.fa���5���P�aǤb鷅����.��[6V���{Yy��ۗ~�p��r��'�"O��z�<���{*����'��Lx�W���I9��Q$�!{:�;̧Є�;U˳ �	���we��/���&�������qN�t��D�Tw>_`��F1�x[ ���bO�LY�wLDh���()q�̨�r�ʭ�3�����$�"���@�H�83[������JE�VaGnW d�2G6�HXz7L��j����SbXhr�hC�Xՙ��xMJ�m���.d����p5E�m.P�/�ub'9�-���o� ��r�H��	9�ޫ~>�dMvE�ޣL��`W���I��%����j�	��E-*�P���Ý���CPMI�~{�y��{����O��?�HG�zǲ�.�o�4� ż���3��l ��i&R�����^���&���R���Ԧ�	
��t���e�x�4֏�KZy��O(���w��ާ]�U��O����s�"#L�v,'la��;U*;;8�%���������OR()E���ę2NX�uNs<5R
�@��-�_�B��r���|'^� ���#mX�Xy]�#9��O��~4�W��[d銂�P~����)T1�"�/u^��=&I�?��:�q��  �p�X�=V��Ν]/(�KU�̈���W�v[C�2݂e���N	4,i��/�Fb���k�DK������xt@�^�p ��9h�/���<3��/����9=�0��sg[�S.�O�I1�B9��=���� �,)� "���ek��[���9���	ǳ��Qu�3���%ɵ�ݦ?��|_Rc�C?)c� �v�r��m��ǵ(\���#wY�G�����*#I�T�����T@���+7�٨=�B��-�<����-�I+80ٕ	xu.��K5���V�8��߮>����N-�zB�+�׸#��0(ޫ7�66��z��X[{U;�c��D�x��p)/<���J�u7p�89�tK��Fr���L��Eh��b�{T�J�#44�~Y-:���(��_(@�~f8s��y���4�7/G�/9W+�&#!V`��U��[���"!��k�u}�@˺'�Iˈ��J&�q8�=��U��������Kk�w��<��}��G��^���9�R!��̢��b��y.�Y���.���ж@����w�t`���T��N���4d��h� �M�@�Yԍ4z�l���ր�D.��+� n��H�M��$۰�;YR&���	.k��,C�H��rVd���3�p�Gu���+�u ;�H?E�TT��vѬ�.x�a0���gɛ�3`�o@�4���`�a�l�0}j|)	;�y��;B��Q�]���AF�RH~���фV.S�[E)�
���X�ߧ�4��y��v=i��C��P����R�P�Q7���o��d\�A=6�)Jɐ�I�;>9�@���;c�ٚ��B^�p^�oƞc��"V�;����WӰ܂���:�}>D>�\ˡ݀�b_��	Ib��R��/蚀�ɨY���(� ���̌x��C/�c�8n�>o�:'��1�WXl@?�Ν$���D�vђ�������cB��m"K N�h�R�+F�� �ݪ��z�&������ 򇳖��k��3��+�����X��x��a��a�� P��~Ye�0L��\�ވ��S��C[*G�_�37�g�t~�@������ĭe7�� ,��FY�(N��$6�y���)�(�?I�J�$m\-�A�r��>�f�լ/`�����8h��+
y�,�z���}At	s`�Ҥ�:@�@�ln��L�����S�ʫ�!���\/�2|D��x��2�!�:c�����*za<jv�X��D������,*s�0=��&�f���H�V�o���̷�q�z �z+�:e����*I>��+����d
����x�WX�
x��W(�\ag��	��Et��ie����%H���F����]�k/���[_�<��/�S�U�	��Jx�曒7�AʩM�
hŤ�хbvF֡S��f$�w5�7��
z}�'��u%�#(�O�qh�$��̆b $�7�0��v���<&_����עh:�a�{�R���9��enb�V��������c�W2jڹ�H'ݕQR]��K[���{Dr�8>2�(q G����jG#@���3ѭO���H��˞й��1tߊ��N;�Rޖ˱���</�{�3��S(��er�mQ!顚mx�yY���NY֍����C�Gǅ�c �c�f���:=R��]b���M�n����"κk����ٙ���
��0���L�M'���]�,xD'Zj�o}�Ÿ�6<�;D���D�7�a��|�,����%A���t��t?}aϭǂu*x� ���#�1��Ss�G��~���BW{
ڗ��?��@S����q�y=�}�md(���`���t�níW�� �Ym����E�mz8Nh_����/j�y�pD��/2/>��x}��l���YI5�|��_��%Y�XlxV64EB    7b19     cd0�:��VT�+星���"�K�P�������4a�������W��Hj�6�4Z�DЕQ��jVz6�G�"�&�唈�9F��Z��,�#�O��Xr�����x _��Ve!Ll�!�k�+iz��&5%�"|����o�K���F`K)�;��F����,����P.�����,��c�~�J�kB�T����'��sq���˕26gh{�ȂRk�&�=ސm��ȉ{���,}����'t�"�����E����tkv�z�����L�����J�yg�ٵ�@�j5D�|dܛ���C��o��qX���)�|w�T����ի�C�V���I� e��I,�nl���?���]���ƞbBb'����&\
Jq�e��7��q�7�}� �޶Mxl�':�������C;�*T� e�����I�A�)�c���?�����)�$�ɺ��R<:��(7�h�P[��5����� ]�'x�t�������֊7��p��&��9����y�|�����޻�g�Q��j�Z�OizS��`<�)��g?p�m���>=�����nG8��g򓧱��Q-/B���t�P9:��CY ���n��3���'��R9`y�p�F�FPp�����;�4g����`�u�3N�Q(� u�TP�-Ø�s�{;���\�Y#_W�qVQ!��%}�
\��E6u0��(���_�������9�%\+�h
���߁�Rx��.L%�Z�9hq� ��-�eOy<$Y-��EA�D`�e9�{�*��)S�#cςEz�c%�5.�h�����ǒ L��xR$%�t`��Q��ue��!k>V�mp���)W�DN����h�a�Gi��_@�5����ޢ� ��r}��Ulh��$��4`�+�x0�����:B�iꁲlzѮ�����:�H�I�,���hD�-�zE��/L��5�UΌ~m,�@wy�*0��e�:�*#� ����/���ƚ0Pl�T0���>I��4"��ù�56�	�u4��kj]^	������fL���U0B��hL4�o2b������<d��B�c�߿�>M+�r)F�[5KP7���ɡL���P �%�o��E�I�el��Һ�[�2qA��.>��`&����D�2�*�y��Mg���c�OQ�m0== �|�!	[��XQ��E7��a�-�>�����-��������T��A����bX��qc�[�1V~�\�X����sX4*�<"��9�8�K�[7��Ҕ��c-h1Y#���_yb�J/��&	W��@N����q1 
/c*��Ö"��`ϰ�d�R�cz�XbAᒄ*/,o6��K�U�|\�ޜ��%X'-��ޥ��D�l���N�Bb0�tDB"~ɰ\�m�v���K������v����� zl*�%/���&.�I:z��b�ww>�p�w���� '|��v{,E��r��"\���q�-Z��G�O�����w!�;4N�L��V��E�ir�H>��(N���5�])��
�T��C��~��_�9���YG��˿�6qg�(�)[�C�Mi�o�@��	-xO7(X��32��ի�u`��BD[��(�Y��n��Ռ�׵����=Д�֤�͕�x�jf����"��z��K5�aȃƄn�nY�����>wo��i�a�5·���52hP*�~@�~n
E9�a27&U%�E�v�Z�6�8���~�����d��rZ�p$��Y!����k�0P�f�v~T%�n�gP6p<M
�D_��d��7��U��9'!��}�Ì�wJ�\�H���ԉN!�`~�պ�TW���^˛�'�O!�p�e�!�kOZ�����Cs�el�Y�Y�J�!Z�cl�HYs�-��%'�mb�4W�=�JA��Z�MB�������zʏ��E*,L�zN��S.�x��� Ui�[�^�'�v��0z���M�ʲI�0=Zi��f����ʗ�������8U���疞���Zc�Q�]�� �%��Pu4�0�L�lJ��8�:{�Րx��J� ӕn���C��$1H��^S��9�]��D��U�~�vR��P�C�p�ȱ���H�售{w����dd`��D6GB����K8
�tZ\ϩ���R���ޯ�İQ��F�`dزL>x ߤ���P� '���[o!wF�,89�	>��}���	�ݦ�
��J���������2�ԩ�v��j���%���c1��6���݋Y>}�&�bH$�c��5z;t��a�D%\,�Wh��+ZU/�kɚ��/����6�˩[�(�Ж���B�M>`��!�=�T���k{2d:�����E�C��cB���1Y����%�%��5�^�ģ0��k��e-���� �c8�\�oh�`��F�7͌��ȫ��U4��Z{s𺫢h|ݷW�������(�\a�Gl��,?F��V�-Tb�X������)�m}c"AM���l(��^&��~����@ȵf!�ԆX���ȳ�U���h,�-�I�?�\�a�Pď��%ɹ�G1�s�D#��Ju+�̺!��
���"�,F��hl��E$�V5��:��^7��։U`��)��Te��0ì]�f����<o�(#)��3��GI����^efI��g[��)��v�����h�c(�J�^ĕ���뫏~��^r:�z�j�:�X � �ea��
��0n�W�4�m��D�#7A�*����C�s����B�#El�X��rA3�3Gd�I�u_  ��0�{Q�5]�MۅQ��ФJx��v�%�\c���I�q��Y�:_'�Q4G,�f�R.	���Uvg�d��⛠ 
�0NqIk��~z�c���ޟ3z@*���Y�gQ�y�GLx{�`�� @���pP��F��#��`�/|E�V��I�� Ua`Lpa3�B�N��nnȝ��Ii�&�;[�;?r�{�?��I��)B�����(��E&�/|�u��u��ΕIps��AL��-�dM�qms7:BsH�\�+��~ ca�d�vK�H��Sy�����h/��R������V|�}&I�l>�d������寡ˋN�DB��'j~���\*��ˊ�,�.��@��˩��
�d�Et�]\��8�P�?ɠ�|L���B��5d��M�͈%P��fF�ƥh�ؽ�5�a;r8u���8ܱ�6�,�3n��}�ٖ�,�,�֨v�̂�,�r%V�4����@l�'