XlxV64EB    2139     ad0�� JS��࿫k<��,���&���cL7���?pc
�p�9o�)	$ѿ!5@�"%�WV�8S�F�ҺY��tY�	�I�0��UU2)o��F3JI�!6 ���y�}x�����q>���W���S���/�7ˁE;_�b#��)��a�=]�ƭ�zg���ւ?����I�J������$������/�Z�jJcru]VO��wC�b0�p�/��6/��(<�z\Qn���}��9�{Oa���l�E!U�w/��+�@����Y����wI��/,�<N����HoəV�ыx�AKL0�H��������|�-�X�e����y�A�^���{RǨG�m�}	;����a,�A���^5�T1����%�`u�����غ�ϔ3	3��ǿ��[k���7Q\�s����b@��C�+�BMn�������:0��4��@��pMAZU@����X�rXN`[uw�-�1q�e���z!6�o��e��Ɋ�� g?������k=b�2�뭺	���M�8j��c 9'�6�g`Y�O0]lL�����dK+ĖO��n����l����Ϡ�@==��|$��@�1c��*u*/�+A�xg�=�ݣ%;�sNT�˺M�]~�J.d��ç�Wj��J�X�� b�=k���B���s@�VkG=N�G (�9BXA5q��}
y�M�4��0��1�pɈ���N|莰r��������{�R��������vZҖϙ�|w��cx9�����XQ�qbVr8KN!�'x��db_�ڷl�`)u��n'K���T�n�����_Y�]:�-2VJ��|�)��|)FqĻ���=�L]Ԋ��v�{�ֳ2�סn�������P��aќ�p��h>p��Q+��l���W$�� �<M��Y��V>I��ތc1&e=������+T�Ԫ9F(���LA��J2�+��i�������Xq����,:<
�%�>`��!�}(�~
%z�b��p�q�fc9�Ӧ>����4%�C[A�x��a�Ra�e�'��O_���&3�{J���xh��b����͸Vu�� &�yBl�;=T�蝡J�=R�������#�n,ȮpD�^k�j�Elh#R����B�kW��B�R������iޛ��x�3��Wp㷵KJn/&TX���2N�Sg���b�n�᫉���h��<�^�h�=b��}�&:45��|�ҚH�q,y+�����,2�6��z!1x���Q37۲�Ù���H��Z�zh��h������$�Z^l�K��,/ҧ�W�`���O���o��	����Ag���7�>��+����5�J:B��4��gk�v+3bh�H]w@�z�Ҍ�5�� i�+Y�|Tl��n������|g�������듈D�T��Vt�,]��f[�� pS)��?����?PT����"$��;��9^��7W����B���/��AsC��H���K��9�fKu��o��|�.�9y��K��.�27�G[�&(f����z�0�bJKV�ŗ����_S&pџR� �_!=(��rIr2w6H���B��	�{HYY^ZH9AȹP�aE)�h"�=ӵ��B�	�۾��Z%�3�c@�َ�T�k����M.�a���	���O�]j����o���\�y����o�r+eP"��G.�\��SW~,�'3���6M@�9Q!���]��k�:|��fVY�;-��}9^����������Z\�Ճiy�b��ɔš&����)�3zD�˸�]��������3�8	��'�i�������_1n#�1�)8yr����nb��F�[��.���Bi<����WL�
y�)��+�Վ=^��C�l��ˉ��UK�=,0�:�悻��|A�M�&Q*�a��:�P�N�	��,P���9���	�ey���W:\�-le��W�ȷr��@�D�m����"+� ��1�!���2�T���;�vǢ�v�=,���n_Ce�|;J��}��F��B2l|g���QW����f���[��x�}��*<��>�)���C"t~vB��~7띴$$�sy�J�����\"���͓v>�G���NF���SFf���0�H���ɭ�@�"��o`ӂ,�����/r.��+�ي%N��׵�<袃0&8l�Ϳ�w@�J�"��p��ߪYE�=o��(�K��WD����Z���Rb(�6ro�-�w��7��؁�������H�V���$��o���0͑�B���A��i� "D��뾁y��([��(���dC�\�X���ZK�'_?��_z��'�q@��I���_�Q���\N��ı�HV ��S�G D_����FDJ�~e� ���E�p������6c�PT�t�v�]��+[y9�>��>x�=ܢ�e<\^��f���v�a�D���	MX(��_���O��~a�.�Ѧv�k��:��������VvT���xhwCg7�R9�i�%�oT9Gj i�X�<�$���ԓTM���qMÁ]!6t��c�'w�%H�?�Q#��ܤ*�]�5?;x��DC���\K�WC�!�����E�F���� G߶V�
�RQ;7^�$��z�G!m�l2��?� {&ӣqL*������ ?ٽ�Ѐ|�A���i�ʹ�/>Ѡ5��E�k�WN
�~���&�U7