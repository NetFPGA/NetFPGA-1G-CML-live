XlxV64EB    fa00    24c0��5���ꋠ>��	2��O�<O�����ˌ6��K��ʅy���$D[���c5E�J���,:� :�1h]c���}_�c(o��ȾE���#�M�;�� ��V�>șL�pC�5t+����Q�3�̾�k����m��%������c~KLS�{�m�-
5���F�<G���{@	-�S�cU���J1鏿��|����&M�P?��ؗ��c�9k�y�5N��v1�V������f�u�|��_���˥�D���qkG����/m�1��I��M�JTa��z�����g ������������Ebo'El�q�'����e�, ^"�������d��6(�U��3�#�J�[d�ɵ3u<` `'��ȧ�"�W~�1�K�(O���v,�*{��V�`���)�$£���6��ǯ�3y �8R�N�[��{��C�1�rDBQ�܁~��mX�D�-�b�7;G����Rқe��y�8S�@�r"0*7 ��1�!n4&�������)�;0��%�fX������K�i��m��g�l����?�K�/�4��	���1�ެ5�� �������2&���\Ê3 kqV�k��l�5�D�C)r�0�����8c֎Mh���yY���J�}��o�Q���ʪ+��
�QSu4�I�xlX+��8F�!L酰o���k�g�q�N	tb�{���k��G�>����1t׀�,��[���6����}���x�3H�;A�y��q��fw�!=^�#�c���d]��Ña��+�5��,k�6o��E�[W{��q�;l�a�!Xծ�C6:�B���F�9�R{|�I/ r�ۅ2�:�R�g�I�����bl�eJl����>doq`��Yb\�����gp�?s��ĝ?�d��'׸qIK8�/cw�^P�)K���F�A�J��82]�V�z���d�Ը�2%D�VI�P���Yq(���R��A�:��ki��s�n3��pD�3���u{� d��~�ځn�����;��X��`��1�g�յ;t�w��kA�˳������,�C1���Ϳ��'����9 �Q�Tnv�_���w�ڀ*�Җ����S>��@DV�y�w�����B���f����f?��S?�|[���Is�'̥�;9���``����#_Y�N��Z-R�&���d�.cSkx2Pp�ȩ����|���Σ}(%����D�-{!�'mJ�����9���>���ۄ��ɒ����Ұ�;_.�m���o|Jjn6�٧��g��U\��Bu'}o�$�Fc�#���	���L�+��,r��g2٤��dp�F�h�m���*��J�lP�85�/� ŽZ�T`^>��������q�����*�5�X���d"��uD�,���"O6���2F��8��)m�F5����Jץ*�:y�<Qe��k�"}m�D1G:ө9��VL�����jb���H������O��$ ��J��2O�\+�����;�nK��T�kQ�q���q���A��7ꉒ5�|�X	�G�/���V�ԟA%e�h�
'
�OC�X��x0*�x�B�����[��hd�T*ٲ����v�=�*����W���t�UPIB�{ <�
��{l�̃�����v��"���Y����E���*����H���M���'�@�:�ݑ�D�c�Y%�����.�}�f��eͮ�,4X�f��|�ϕ��]�n(��s��ǅ�V�;�t��N����,G<m�.XQ�V`��w�w�k���l���g�si�
�M���ߺ�Z	�����:f"�`�ߵ�k�<�dR�Xx�wR	�i �u�n�N(O^z��{/h�
#O��#�
� l=n�\���n�m��m����Tn����+����
D�\՚^�i����C4��K��;B/�����5kS	�,;s�	�)���Gf�MB���E#4����Di%���)���96i/����l���("��h��i]?���m�ύ,*�Wem6ܥ�Y0������!t�8�TT��E��U�4�3�� m���|��&���}��}����F%��w\�MM�SY����8��� fp�'��m�r��+����o��7�ę��L�׌g���G	��\�V`�ں��E���K�tKCmob���nDؔM���d��~��w�]I@}��ѰB��D"�������Ơ���㧆X��$�����:��XV�O5&bohv[Kb��sc�i�+�C��4;<���&��'�4�%���c�!�>'���v��S�k�[������6����b��I��0���lq�bmuO���xa!e���\~���-�f���h(�&�^�-G	#ر�u-��z��C��>�a����5���_�(q�_%2��@�<W`O��(١���i\���_,-�g�j?���"����J ��}�p���9�Җ�{ �.�YY�!�|6�!Ne��;����H($4�!��V+502|��sڇOc���:Y]n/���"K�&ɻpW<���@KN�W��"�j��k�ZW-�3� b���Dz�ۖj�>��)V�}�Z�D��E/���u�?!�Zj9A{;���^�~Na^�ְ1�=�n�@�/

nݐ�QB�\ĎQF&���;��x��;�R�]f�j���.f�U���q)��>��3锠��GYo/�6m��s��g���6�wE�v:E7Nw�P]]�1��mO��jWo��[���Ӽ$,��#�k�:d��G�W�`��GB>�h�Hk������q�xO�yh�#���R�Mg 3�͋Ϲ�r�
~ؑ���m�MM1Qӫ�E� �H�+kyd�q�t��������+Ih#��fQ4����ҷ/�fj�Y��	�����T����0Y��8+kXxW�=�l	�y����?�D�3Vv)�}-��퇨LE�=-.�e��Jȹ"���r��T�JCz��JRh��(u�G�#�فދ��I"iм�����F�$Y�ƿ�@_��*:"5����1"Jb�e?���߫���;��-$�Ҷ3���DOZR�_��W�ޢ������UC{H=�m��
�8����?$��EBR��Ѣ�W^�l�i�>�hr���Ǒ���`p ��%F��
\���
_R��Y�x�QW�p��ϖ��
�l���� 3'���_��y=��JVǄ7�3ON&�~	�]l�Ӌ�1�R{�@�D�bR�S��g��#��'>L#AIoZ��S�w�vܐ��N����E������&鈺d��ϗ�DE_ܳBC�w,Ǥ-p\�8�ʪ�ڙ&6rŨ��
ܠ�U#��_����%�A ��H�R8/K�p@��M?�0Ù�D	���O�C;�����W������0���h3A�7���U��B�FO3�����d���ƭ~_�Z�N�)���#��v�Ѭq����~��P���s�#�����N�<ë#�5�񰄞�NGY�WFfΏ�zI�><�%���Yl����k��\��LL� �Կa�̒Yja�^R-�9�ld5�歽Q�a�,�÷�Iu�Z�KD��C(�feǪ@�¨~���{��8�'!���S4]�*�7*�s�mS+�3qM�(7ʧ�E_7g�H·�W�ƈ�m_s�]*&V�@k`3x�;\0�%���c�A��rǄQ� �{����i����(�{��ŔoD�R~CӎcGQ���X>�0|�%� ��]����F}��������a�	�d�� ����OF���E`m�Ym�������j�Y��凱qPRV䁰��į���bnX�� ���2jN7x�_���u UoFL�Bw:�®�J��"��#��Z��L�"[����Y�Je�[�*𙈳��^ڑX�H3�5,-�Yu]���������������j&��3T���^���e~̾Op=�����[ہL��jL2j��?��%��{��'�!�[4���w�� c��wz�D]*jA�JoC��k�p�XU�{�y���qtD�j��rf�!Pny�!�i�5�V���Z$�����6���c� �c�P�_K�]H�q�]��+�_��c@�!F��qH�czy��H͖҅Hp�6i�nu��ɯ��U'_aӹ_Ͼ�O��,^�N���֯	��`��_ױ�f}0��Ȑ�y������5�yxK�Kb�M�H��bҠ/+��,~�j��]��0�wzh���Ԣ%놕l}K�x�L ���6����.��!��JI�AQ��˒ۯ�3٨)r��Nt�О]��o=h���/�Z-�gOd��/�NB+Z�@$�35��A����s��	lݟ{P��I�{���%\C3�3�m�@�jj���'M�+e��ӜK@����[��AxbЯvT�V��/���_�����UmXt�t�v~���6��@����"�C<>��V��
7���)Ȫ�F�f���@ta�Ys�!N��ߧM�4�:�u��J��@(=�,���
�UM49 ��Ē���t���X �&x쏶}���l�敋�Θ�F���7��L�"���ʹ�f��1kF��;��`k����N�S�"��$�u�n�"�g�ĉYS��ݝ3}➽l;�	���_��z2E$���*�Y� ]���20�� �E�P�,�fn�qY��6���W��C��i~ŻP�u\� I0��?JĲ�4Y$A?�.��7��.'�=���PKAL�L������\n{ ���vq�����?_5��r*�PA ��h�D!�JF�]1���5�[���@p�Cit�X���T�V�����m}���lº/��帞#n��8Z�,��-�	�f���F0��
�Q$��o�t^��Q�B�(���]Ye*����uk��!s���\�t��c2�4�uGf	�T2�=Tȯ��U�R�7� B�����GOP\N/|�v�E�K��T�D�TD����2W嘤�}�`X���yϱT)�~]�[� l<�V����s�ehE3 %WX��-��<�m|3��d�VU_���] a͠	a������u%����r;��_�B�G��WÏ�'���8%��7�l(	�4��p�����,�.q�qk�Ih��W@r�]��J��y��p�ե	���b�K*��cH��a�a��������Q��Ĉ��=Q�u߳�	{���~����.��LW�Z�_���3�,P�Q�>�����9�DwSF�./H@���6b7E�Z�fI�m��i�E S�5x�	��>2�Q�>���=_B�\韅����b?|vӮC[6��<�`Wn*�n��C=+�;��sf��7F�P�P���>�{��
�BM���x�K[ϧ���a�%��HD.�
�:ߨy�ǔ~���O�hR�르?7t'ւHn:��]D�4�`��~����Î����f��_g���M���RH�|�҅b���X>#cn�W%����pZK�/�_uB/�ͳ驳mQ�;3�DSxb��1�~S�Tz]Y�L3DF��^�f�qF�;��&�"oZG�Q�UO�$��!ξ,D�c��}n�#ׁu6в�,	����+\:����B���C����|:��mw�E	ĵG�?��g�&�gg���1�]X�g��~�{%���[��r�<��@H�� �D���`��E� �q�٥U�i���DT�/X���s���u�ޒ:�:���/�4VïZ������2��K7��k��Luc*��K��=R/8kYvoS(�dC��$E2�qoßڌ8m�Q�=b*�Tx��ƠOu������}�H�W��Zw
#��"4M���7�˕e{�E������NO��䬔[�������+�U���iך2�-�`�C����>N�?G�c�t1o�O�R����������q����/�XH����C�`���iR괢�[��J�=N%�yJ�������� "6���d�M���L�����#��3�d`��b4yT�֗Hv��2Q�0�kk�🯶9b}>hP�q�_�$(���=1�S��������BY#M�A	1���pI�o��a�G-��A!,�,Q���	���y�O���B���SW��������<�(͎�\���У�`y�����˰���X�V玩���ۦ�C+�����j3�{.��a����L~��D��X��_)S��	���1*�gP�'���/%��B�(穆�nym28������˥~���ƥ|0�o��X�^b�	�V��F��T��`#{�AP�E�
��t�p.�N�O?`�}S�S�����!�vSs�M���)��A��L"?�*[�~�W^�	k�5#�5���הV��C���p��?"!����"胼z���p�F�������s��|P��~��v�L<c<
����IMe=�ILm��}(�k,z���B�-Iy���s�2�{�0�j⻒0<�P��w;���/C�FY@7(�6�;�`��
�!�I)����'w�j������������d��a�m��!�B�� �;�̪Kzq�� ��@q�l�F&����t�R�D��+4~H����������R��>��r�4B7�O�5̌���@Sڵ�<�a93�+�u%ѿ�P�I����Jݱ�1�'ԭ��5hb)�Q&�Dy����?q�G�4Vܿnj͹�����&��ֳ�{��oUZ7X�5 ��t�1�����3�<"݃�֬�RS�l�[��#��f� rN�	��������b�pͼ�y8Nv����K�[�᎖W��EiC�֣�A�'Hd:��A�����ߚz��.8��aǢ�r^���?e�
C�9K�w11�U j�dl��j�Dҫ60���n��h@X荻��M>������"���%�F5��u�s�p�涄nC�2җX�kb�V1�>���$/�e�RO�p�j��^�IC��TQ�	L�}s�����#\��.��%�n��β���.)[�th�b�բ)��G�Sa���"  =h2,���I��۩	�^ը��~"%��$��q������'[����^��4��_ק�n��@���+m��_f�d���|*;�]*^����M�����ݒ _6"�es�ȁ�����z6�\"�Kb2�P��� �0���]���	./��[�]�=��ʀ&�g����83vl��4���˫�h��7M�"���]��Ӵg��	e�a�T�E�3f44���֚:��l%�=�'YA�����U	�dy�w�$5����[��vN1':�$�*��g���o��PuR �^1>�1\D�@v9�(a1]2�ć�!{O��ym�vi��ɻ�ri��b�����m�E~�D��vfZU7�z-Y_P�Rf�P������.�GK�b��"1m8f��I[�%�9�F��4�j�Xcs��U�pP�H^9f`h� fbٌ0��-Sr�J�<HѮ�1f��� ��|H�Rb�]Q�;�J�!��I8ol�ۂK0N�}�����Ʈ�6Ѵ��>cQ
��e37,��`��*��JC���᭍��@�v_�H!���P/.������W�	�'U�}Y'�l������b�vB������hY���X�d��?ڨ��������'C;�f�CNb�C[+t�$��c%��^����P�PSj��� ����:r��BiG�����wA�%����P�m�7��B�Z�tʾ\d@{x����c�$y�� �I�Ep���J�;��Y��%v�"ݜ{�7.��:�q���L;e�����l�zW���ƈ�\;ś���f�4�f���	l=�)u��]J(����O�$��E��%	kT_��p�k9���(I��ܟ�q���ҍw�L�_�-�	����se�����Wqg�1��]�l$#�t�`��R0q|8Ad>��&+F�*�<�WGo��K�D����m���%5��W�y�k۠+��I)I���dO�F�JqoM���M�HV�0X�p556��$��7=fG�H@�ֶ]ʂ�>eX��zG�,��庇_�+�m�`A��>C�4�'�KpyG��q=�p���S�CU"��m��6Ԓ�9.�	����]��;+�^O��!<8��W���7n_�W���j),^�x�"W�#>f�#���dO\�Y��mT
�S�-�N�2q�C�5�Ƌ�J�_Y�|p��;�>�<P�A�;������nk� �u)x�BD��VY5PS����t��	|��j,M�v�x5��"-.��4N�HUdO�����C%3�O�窯	�M؅԰����73@�s�J�����3|�7��U_�N�'3 �>���x���j�sZ7��}�Z�p�g#�����ȱ��j�zZ�n(����Q�'�\�F�*G�ZŚ�cЖzrx�廐RO�:X!�H�-K�6��Ŕ�:�*zO>ХD��㫴� �\l�zr�TAT����Ύ��]yry�9��^��=c⯴���\�$�?� U�ճ����b���oRs� '=�Շ��X*ݯ�Ń���|�i�8F��u�6��e��Q�(]0�c���:�~J����I�#��}3�jC.�{��סt㏥�q�C��f�H���d9�����,��t�N�K?����`la��Qi��X�����aR<�����Si��eo)6[�k˒6��R��ݷ��a�⾯��Z,���D�KE��|�����Do��o�Ţ�����!!�u�}5��y����B��Y��z{q��D[壱n�V�Z���1�z纾����d�\q=�� �'�:}�X "q���^,�g_q� QΔ&���lQ�������4�`q�!�&�fY��[P�q࿆o)��Hz(X�/����C�M_�w�/�<�+f떸zVٵý(S�\�	���G��+gu�"�7DR��E�V��D>�1���+V�+h�.�\�T�.�Ig��ѧN���%=  �=[���W�$�f��}��U@�. �K9J\Л�f¢��	JiyhT,�~5A�r���y[�~�~  E>�X3�
0�s���+� �f�/�u,U�tƿ2���	�RG�=�yu9�ݸhW��VZ���	ґ��\���D��ZCܑV�*�����gRO��.T$�F�Ќ�;H��r�x���ʖ���Ά��ԗ��+-���z�غ#���M�=k��<%SPF���PE�:���.�wHW#���DE��-��v �"�./��Kd�'Nh����V�u�UsAJ;q�L\��ɵ�`(+��ʊY�V+@v�^	*�Q~��^+�j�͢܄���0x�n���XlxV64EB    fa00    25b057Ƌ9{EGR��d�%�AÁ�����vη�h�3�����C�J�A��5��7�w$71�n��&D[��̎d�7��D|)l�y����Z�S�+�t�h.�gp�+0j��[F�f�+������4b}����~Hq��~��a�����խ=݊�U��wm�N �T�	���(3����iS���K� ��FAR�"av���f4����GE(d~t��N_�@〞'���8%+d_N��~>��68�.G%R�/`#���ߏ0h��>x�[�̩�4�k,?����	��2�����m��3)HC�}��Ы��9�28v��'/Bϳ~n>�c�Mg���B�#�q�}��ڊs��+�R�%����	�DE�@p_��b(���Q�RIf*2j��O��4@b��v�;B���k�e��r,(d/Q`�a�e���MI),u^G���B�ɣH�qe�7vľ�n���(�ei�l����GtC�:�:��:�P��[B��Kh�m��h��2�3��Z��ߠW-�:�/������/�[�G��(sdY��QR�<��q���7[��	��a9!<o;���I񺲲��iQ�J:;3��a9�s�F��lk�E��g6�s��������pS��>(Ҫ�<��e�l�;�J�)x�����m��53v��A�k8ZTrJa��H���r��m\
OǭE�*o+8oǂ��:�j�j����w�{�g>i�8��JJBN??PO|�����~NZL��e�W��I�E��Ȕ���uْ��IOP)dʂމF�|�>>p������g6�F��Q�b&������;��zv�;xEP�j�I��؏��������U}L��Q�
�0�&���h����4�����y���$����h����f��Ot�n���H��=�$��#�������@�]���.��!xHAք���&��a����ע����v"Ϥ	k��d����̷ ���ϧ��t�}�Y�5�����z� ���hs��n��5Y>�&��GUP�#�0cz� ݶK2,�
�m2��n�1� Iü�-��c��+�/#	Vh�^��.5�z�ȴ���;	w)
������b�0�[�B�@0��?4H�oi��k�X�r���Ԫ|�\�>�֋y��FeX�vT�/Q�1�{�D�GbåW@ba�U� KLU$*�
(&����¹���,OO�H4,�Ks9��~��S�}�\�$Qҏ���m��A�Sߺ:�7Q��#\���z�q T$_�Ə&�I�}W [^��:r�j������jt�j�9�z���!��!>[�weЫnE��d�h�9��������I �
��WI[t�~^A���7 Ш1��ﮍ�`������J�O%�}���DHRjT�.��iU�@��`�'�W/#���J}�N$|RVů��|�׷`i��`�ar-�<��j�ڋ72?!L�2~O~��ը�Sy�-Hf�J�5�$�p�8��4��l��P��{��z���fਙ��dC���elڵYO���Y��J�Y�$�V�ПlK2���9�8j�.�-C�tv֘��¿tz|wB���
b��p�:��P�$?2���5-� (�>o��*�@C0�Sv��O�Y3��Y5��DA��"����@?p{6��r��
j��|�}Au��~]"�4:���!�ٵ� �����K�[�2�o�K�`#W"�z��B54�ȗ�y�g����E(�UR+n�*��s���=����4x%s���T���	���h'L���6�v�?m��i�"��
<[� ��d`���ݟ�[2+)��&}�\��^0��^�:���R5ˮ�"JDgGq��>�i���ǑM��C��A]NVȂҳEn������]�Ȑ9�I�����R�M�b�µ2So$�=?��$;���P� N��p L�$�wJ�{���`y?R^ث:v"S�j���wD�s�&�Ǜ���p�1�� ��[��Rݴ�P	������ξ�
�Bw_.�[�1�4��V�� yE#8�}�OЄ������x�6i� �.�hv���M#�Ȑ�e�*H�cZ��Q�Ԭx ��W ��!�G�7�<��E���'g.��k��	����� �`�_C�3���X���RIf����qz�^1��A�Z���qs[H,�!jn^0�y�b9t?Ȓ}*܆�k�߹�q@=����L�p�N}�,��������������Ļ��
�ѷ��	НZ�w��Tk��z�m��:)�
�:���ձ����Y��|�kI������$�P!�ߎ�ƺ��&8Jt?��P�9�_��S�˗��Fu���3���O�8���5��eG�@�e�^,b��� �G�Y!�ǽN}��c4��B �y��s��3��W|�LSC�u��Tp��oI��O%�{;T���	Jqћ��K��>�������hFv!�@�,ö%�bB|�dx
��t;Gя��]��~%��	i8�cᥬQ8ٚ���Ue��Z�Lx��$��V+0�nb��}w� ~9-�J�":)�QN>�����P3�����t�쥛?y��L�'��(��_��Ajl7P\k�40��<�����TK�z��'Xk\�4��If

��u�k:�g?8xgc^'f.�t��u_��v��E�4K(���E�>���=�&��	��Yp�;f����� Et9^s�Q�5@�n�$ш��8�������f����̞���#���텴^�=z*�s(/���%�(J��f�"3 �'W���4��.Nݏ�WKd��)rl*�^{P
Cw�Μ�X4Hp=��ρ��"Gs=w��o�'[~ F:N[�6�Z�y}�4yϝ���Wu����hʴ��-����r����6���5�
�}��^��t���s3����;�?J%s)F�\��{?=dmJ��$��|��\m���6r��[�PІ˩Y՗Z���	�|8�#�~a-4�}�i��xӚ�ސ��l��Y{Q��� ry	�<zf�{W9ܫ�(]R>�9Hf�|�ysZ�5��#�"e<��%�#?�h�騇���oQ����l> S��w���X�Ȍ(��4Q��G�q�d�����{x��l�w
`bm�a�vw�Y쓖8Ń�e��rj;a�k��1��~������u����Y�X��7�|[Û�ܱA$����BQ$���Lg�������w� �N���W���(�3᝿��'��x'T۽L`f�����t7<�����50�+@���`������>��>��T�����9�@v�C��r�Z-�M����P����zl��ɮUU?���|xk��+��	�ix�u��F:�e⮞� pt�>�:�q� �VL4�H�ǰ:Ok@T� ��+�
��n�bNڿ?	�����dw&�JE0u��=�(�JO�hqiKCߎ��O�k�*4m0��d�3�j3*�i����MD�N��c(�ͦ`\�;>Τu�UHZY�y��S��n�����/#$)X�&�Ώ�=��f�qd܊��Z���ե�}���h|�-��e�mr̸����3kVm�ۀ$��]j��s���[�E���Ή����w������/	�h0�t�c�bA��W��j�-�f5�XU�Xc7��h��*�q�^!�sU6�h�|�������މ�^A%��4�V�|�/�`Ʒ�*���Uy^ ���_h��~�����f��h�������4�&z����8"��\/?�����;�~ٮ7��>l�Du8��	<f����v�dtG*��X
a���Ӝ���u�_
A>",D��4�Jp��{j%+��ǵt=���~x�8q�#�T�J8�/��ρ��00E�����DA� �]𡫜����B}WE�YhΉ23�e4��|FĦ��V3��/I��Ի���N����'[�j ����R������(�I�ǂ4hdk%t쁦a��ms�u����>VX$���M2��l��Z���[]�����	�g9~��\�a���T�S�	��$ﾣs�x���uQ��3ؕf�V��{[|�G��Ά`r��o�}��Ӝ�i~qʇp��u����+9v��_��	6��G���� �\>2�����C���@>3�5��߭.�6{0�
�G-������\QQ��1�~m��( :�j��~�\�҂'�*�1�=_t�V�����ʒ'褫��fEk4�E��[���34�̌Fb �|DBhW�̍/� �Т9��̭*C����2���]���tqf�?B0��U��ݶ�Wg�I����1����[|H�t����؟��"�1�Π�bbqC�ֈ1�$�"���°��%��������>���hVPV���j�?���O���8���Z|�?��Otk�,꺇a�Xrf�̤2,m��ߗ�i~��s�ۈ!-��l� &=����k�]W�Rq�)�q�ݎđ���eѸ�iM��?< �.�e'�|� ۋ`ʔY������VCV1���\�����{�Y�2�+E[�o����ľ�+23�$�!w_��Z��Ǡ9����Z^('v�-�\��
Jk�Z��ˏ�-u�4���b_��v�����0�O��u��N�BY�M@R�N���z����2��@��� �Y1��N�Y�-qt�]��(��*ZH��nԨ��})��W~N�9??ux�q��D��i����a8<<,
/�s˘�������+���?l~�J�-v2��ߔ����Q M�\C��r��斉���Z�ʇP�m����"�G��+��y�RS��� �#E�H��	sDz7]`���W�p3w��%,&�-[�?�M\�n��T���ê_;�P���eT|��8�e�J/���9>#7�lY�{*�qoZJv�~��c�t�k�̥UݙTE���v�`5���e���R0���ٰ�3A	$�����v�*�o$޳t5S��nk�7��J	��t�3�`��+�D�J�&�{���<\��o�w����ҐQ3�9�pG;���s>���j� ѕ ���}�\��jp���t���M���'5�6�.��c%����c/$e]�7�x���o>�x�`O��0E�����|�𼒵��rb���-;���x�d~j�T��Y�L�^�2�	,-�ϯ��v3~���CF��m�:_ғ�A��j']�l~܉�k8��&��uO� ��_j'����.	��R�`���m�"ǖ��a{+���Dжu^�+Kp1����,1>�9���Br�p(u�a�W���ڻmT�b��Yx�����/�@�</�`��k�黒6��	ki��5㹏�R���Ow�-�����b�$+�'�=yaw&�^��,��'�/�y*z?ܵ�߉�����Ng?T�PR�.���Ǻ��`J� �t�b��U�ne��"��v�����*�U�j@����	����!�cA���
l\���6��"�(���ܬc�`� 0^6y9mOFB���D�g���2T6r������c.ǝ�Gj��.�)���-iI�0J`�:��m����k�+![�غز���G}�,�G�����	j�v8'�[�=��}�]���'#���˯!�r�e/�dXxd�`���ws��h	z��(\&ZmQ�w�b��N<	���U~Y�U#���=9W���0�K�.8���FZ�)o'6D����S����̳D<rM��y�z������c��p� %AԹ���������q�R��`up����c53[��~�������'v:�����9�L�#M;�(�(���Jc��
��x����t���b�[O�^�e�;^�5bg�r4Z�e���_��&��X������5�%|�KW�"�n�&�D�F�ʽ�%����Ҿ�2 �SC��C��)������c9[�.�~�L�� (��?�,}�w+�!�!��LW�E����t�=�Y��������w��NGLK<>2��:����F�e��9\I�����lh����"������8�������+?�
v"�Q�� @���y��$��9 _��a��s�x?�����O��{��Y�(��|\�`�? zH� �$����]���jy��&Oẗ́q�G�OD�8�;ņ`+fCL�D�Eӟ���Q� 8A%ɵ	��y��=���������0|�����H7ks�b	�R�c��<$v[�A\�7�����Q`�}��%B�A���K�n�_O���.hi�?w�Zu�m�&�<��*�O۝Bi�b+����ɗ`�4��L)m�kQ���ԁC/bqBW��`t$+��}Z�ţ+���9��M����T�Q�5I�T��E���*a��q8^�'Ei�6s!_5Cۍl�TO56��~�8N|T�	�fIq{Q�>��w��3��$����I���s��P��q�?��\��-K�&0>p�������8���Z��
>��8E�+�7n�r�����t(ǒ	9��*y��}MI������~�Qou�T ��)�%7�ϖ�����(dxE�_M�W���KM���|��'L;0t;_᭜j�(�^�Ffnj��zx����.�N�΄I��~���bJi�� Ի4��l"����
�U=�����ɯNgb�0'�i'趰��Mn�HR�����(mG��(�nIR"���j(#�=�q�f�诶ӌ�Z�͌�`�'?�'=i��*�v�@�res'8��~P�7����[�KgB��~w'%�L(K�{�����H{_�(͆%%�!N��8��KiX&�C�ou��(��Z<x݀%M�;�A���Ǭ��c<d��Jt}zo����dV�l�!B��&F�QF��틑�B�=T �؁z���{�ޤO�A�|�Zjs�O!	Y_-n��ea�����0B��F���~�W ԥ�������i.rv����[�7lJbB�ȑ�Lդ�\���A:Ie뾽�!��#�.����5� (�v6��/���'�iݿV 'Z@�ǃ�}4&q�X�BQ�Hr��_��a��X;R������wlog�>���#���A�@ޮD�+�A!�'��eL���Z�u�,��)$���cŬ�V;�\;�ZƎ�=�5�rhG�x�s���to�1#�MT��S3 9S�_Y�ٺ��:������M9pwt¿������[����BM���v�B���r��X�^��6�j�hR�[�x�Ӹk�:wz��:�������x�E$�-N��dj=X�y��8 G�����
�ĭ�~���k;lk�n�eA�_��!��d��G�ő7H�o������y�����!9B��ӣt�S"<��);y*�����A���S�W�L����w�[��Kh�ϲ�+Kz��߽n�{Z羁*���I�]��y$T�����ZB���rd��e��u����	#� yk���<l[�5�17aM\%�b��YyA�;~��;�ݙ�͐�<[!�O|�e�zb<��F��X�T2	�J=�DA~	�nl2�;���:����m�o��A���a�����mQ�F�\t[ҙ��Ya��}��X�����|O�Z.XY�x����{v_b�J�N��p����hF���zxF�v��\�9v�k�=�����h�"��'�S^�d,qC���`0	�w����G_��E������'����k� �+��;�֖#�DE��R\��ObQ�_bM{�za�2�@+S@��7�6�wT�"ջuR��߻�0Q�Ck�eq�W�d>�-*��~������V�I�ͅl@v�H�B�,
�:慨��YO�������CW�<��{7.��z��B
�'�%��gK��
�	�؝\�At���6+��f���Z������3Fk���~H6	nzDf���sJu��CeC]Nz�"rj�O&}����r�3�� e�9t�{��N
�9�S�e�H�	^!���&s-�U;@	2վ�RS��.9�"|�&a�q.H��}����u٧����ƋV#�냲2���.�\����5@���ǔ��=�G�=��eq�Y�{NI����Lh慎��=Pu��H��w-&�_�-��թj�_�uk0���L���w/�%U8�\2���Gg�YKA.�V��(��k�m�?f�A̪�y���b�0����խݦw>�d�AL�&�G�#ך|����q}�̿���5��~|� r������e� <ӆ?�*$#i�ѣ�q+��F���/g�]�	L��y�R�oc����$�u_θ��6=
�,�.,Q�qD�װ>#(�ε9?V�����xP:��F�WE=ϻK���� ۩��CJ�!��<�zu���7��`M��V��q�":�W<�;J1�c$$4�Z��PQ��������c>D�)R�ĈXz	���xet�H͞�;�����oTW\�*M���U��[�V�uף.L}�&&�O`d�v�4#D���'C���$xbᇯ��~�i���i���	X)�����{>v����)��g>�+�e��/:3�s�ݘ89���,�e�@4&�C$CF,σ�X*X���w�nl�L؟�N�U�UVP�Fv@�qʐ�gb/��^����D$"^��ؚ�m
r�]�Y��]���!<���D����Z��9�?t��t������`6;��K���!��t��қ�30�sj�c����f�Ӗ�c�'��U}��c���1DD���b����	Sg�g�)�TH�'�oī&�0��5��S�Q@/�Qv��7zI�+���6Y�+@�4:gz�X��   ����J6��0h��VmF�0L�p�?r%���W;�Tz4��9�k����W
�ee��GN)e�C�
LsJ�������A܍��X�{.�o��J��9������=��G�5���i��Y�e^����7���tx{�aw�3}.�Om?���8B�M�E�5'��'�)��J͆o�n<I$�|�"��R��G�7}5z�t�o�	�=C�Jߏy�-<A�ʣ�g�|ߒl�3~5�y�r-ϟ��c�����c�e��y&�No�p �o��I��јx���Z\�/ga��i��Y��O<6_o�3IH�.1�]���ּq�%�@s�e���I7��6����a��M�d!��!�)�މ�
{E�5��eiJ��S7ճ}0�<�I��~a�`Ygo� m�X �/��kR� ��+NY����!j��A�
=1�m�]]�@7���&{Yt���N�ipR�����Uv���J��� ژGb�ɔ(=n.��b_�q�7�O-]��:z�۞7�!#�b���[N��ȓ1�Z�ō<i���_"vi�~�&�H�[�Ֆ�B�w:QCԐ� ��\)jY��K,q�MU���O�R�|��ƈ��޿�ފC����0������*!3c8���8C{�ɏu5xo8�g����|���xv۷�y5v�(�@"K��@Yٕ0?�X���x���i�A1���V��tJԵZ\��1{~ p}�ѵ���/���:�RB�Fd����Z�'�)��D��ՑwXlxV64EB    fa00    20a0�u��n��w������I�Ё>x��'�>|��h�b�29��7�܊�^s���un<��q�y����5�R�ήYK4��3���7(� �Ց�V����g��bbR�1pY����� ���V%g�ps0���	?[f+y��n�VD��ڦhe�M���@���^���ABr���ش?��&t�?��{�x��b����c2*J�ߜ�.�e99p��L:3OԛP�J�&Ä�$뜇�#��xf����V7�_��HL��뼋�x�Y�E>1/[>���b�u�߭,K���
�l�R���٥0�x���m87�{�yt��gg�����A��@h���yXg�/n.�1W5��_�8�.�����gD#񂤽��h̲�**�{�ǭ.V_x/ Ac�zЭ��X�zٶ�}�,����E%^{wҸ�8Q�4u����I[�`��q@S���e��I��(QU���Y�`�r���oU�)�z}5b�G��֘��yR�?k������-镠'���]W��0��_30�P�N/�I�h:=N��;/��3�J+�|on[�C�Ծ<C��HZ��}�XF@}ss�������xȬ"��M̓g�09�dL��ߨ��T��۵�U�� >2Cf�
���ZP�N;Vo�Z����.3_��ʊ�V�2Gf���ڗr|E@=�Ћ�^�5�sJ�x_��{��O �'L�i�v�D
>��O����e�S���6���FW>W�yP�R�B4� Gq����D�&i�F�S=5ٛ��55��l���n�R¤����З�]���]�&2�9���^48�z�͓�UB�W��&ʕ#a3��fe[ �=����12��}���w��Ϻ�e`	.��NŌ6@ç�{�N� �j��F��q�N� ���@�ZP��6�nfrY?E��K�K�z��OƥFI*]�L$=nਂ�7��᳟4T����o�e�=/���VԺ�u.0;D����6w%E2�Ѓ�}0���8���)XZ��y�7.��N-���ȋ`�i��ף���O�7l�o�����:��$��̔��L3�ث܎�����/r>d�֪�k`U���Kzk���Ɉh�	���H���N�D��	�e��l����`k�;qj��d����Sj�V���kS�1�1��6����[o3L��2��Zl�ΪN�ܬ��Y]l�[�l�ܭ�d��ՂO4Q 2��[����V�������?���J~mB����\��w�Sz���tۏQ����7x(T)��y�I��Y��-�|B�=�38Ί��aW,@�ȡ�;꿢�u�VC6���[��o�Q�z��=N`gr���O}�{���xF`�:�ΏU�h�������%��[���"-��0촍������Cn��mA�aW��<)��bZ��jE�+q�ճ�JhE���_ 痋.P�	0��1 ��a��oV��M�{o�8�$�,?��|r�>��O�J�o<�k9ơ���]m��(��7�țww�;&N3�s㐕-Y��5;\ӏ��'��U!e:��`����f6ę����/b�� �Q��Uܿ��6�n�\Hoߑ$w2@t�O�ݯ�0?7��*IRK9I��$��e�I2�NeR�S���-���K��I�5�@�D�O����]�<�t�z}�Q6&�%��%�T&l��<��HO2����w81Ť�_g��-����:$��e�QD��g�69~H'Pg�I��:� Ȭ�؅�����9,�tgP���)ڠo�%�xkѠO�+
���(�p	�	^�
vCWip�~g�:!�D 	r��f�E�����
����ゆ��\`S& �Ε���.�"!yekeRA�t����T����e"]��v�Ww���=J.'�*�p��&�"�~�~zp2�Q���"�,�[�������F�&s�QB����yC��a���ƙ�3X���%m�5��j�r�1	v31��%|�w]��</X��U{i�{��N����÷\\���/�N���0m �����*���n\�
��Ǿ��1n�*�l�0ɐ "��U����n�Z֕�x�J-�Ϡ(
$v͐&��`����ጥ=���E�i�Z}ڜ>�#��tn��Vm���*�$A��Ć/��c�ا�n��2
����BxD��yL����W�/��2ɟ%�a^W6���(顦-��Ht���?�}����ߌ~���cۍu�b�"�2� �4 ��}F�%e��'^��O'o�)� ��E/zeԞ{��K��Ce۽}�;�ýk��xF��z�@:��rpH�H�s9_���o/�P��i��c:dTӨX+��-K�^8{�3�~a���ӏ�@�F�A�^�I&�.%Wf�a�R��|G|�ǪJ�΍�}P������|g�DVA�iCǯBx�����x1�]�L:�]E��6:<�g��/"���eR��7m��5/J�����#sw�˛`X��q0yL���dHxJ�;4"z��˴��`��C����l�����٘m�	�_� �[`g��se�����@"TD,����n8�~\�n�)Fe�Ձ�/#����T#�O��fD��s��E���Gg����ob���.H�h�?*�k�)}�M���,%��"��o?F|��p��ܽ�B�[0	����RX���T�ɳXv�6��V<W\Ӑ��KxO�����7b�m�I.�� W���r��[48��+�2��������� /5ٔ�n���gj`s�����M�����oݝά�8�(�@�5f�8�H�����Δ#R���IH�RIH�^n�m5�Slݱ��&� �H�{�-��"����7���4�?U�/�8�+�U��)��8�� UD���������,��u��M��Uo��u��,�j�ٜ�V3��+�0�!�!"��j��%2&r����p�q�㧼'.?�6���^G1�ـ�^�F2m� F7�9�3�ȥ�4��5�FM���;9	ȂDiˮC/s���m%@�7߰�U׊T���鉙���wE�˝�_�I�1ᡬ3�~��~�k��h�>YF��f"H&�� �+	��*�Qbͼ,
�M��b0$3�5��ԞDKn1����45p����Nt��qw�M����u�Ф�j�@�q.��
R���*:+T7�YG3��&?�af�Ԕ�kF�����&@�B�#���I��
\R�'�
�R]vy�=�KZ�Cn�ai�	�rpQ���E��3Jt>{�MD-"� �%B�E�H�	Ed
ݡ�6`?|��YC�N49X���1$���T��~��'o��W� f̃NDJ��
�E<ҏJ�?�s8唎��E�h[`���2��D�	��j�x���hG�Yk��[NxRdR!HC[�PSZ#�d{����<e�~�<�%�Mzj�LG)X���r���T��7�k_9���uNN����e�s�m��"�0�Rd
ͫ��!8��It��zr�,G���v-��Q͵��E��E
?k,UC�x0���L���1��	Z�=L�o@C�5�\T{��:��V�}+�����bm��RF� E��Zq�M~q_���Ch�5��sƕA�#�,�E�l:\��*�"���Z�ҭ�X��J�(�S�קǛFt�č����D"-���g��w��L�����`�Pc .��13���-�R�@�Մ�9`������8��W�"õFF�bV��Y��3o�e�3콾�ڤ2ř�e�;!56���%_-G����j����hZ�����h��m�h�E<�e��;G����DQ5E�-$�z^k�º���M����g[���t[��$��Q���r�}�^��F�f�Q_�MV�3O2'e�z	�\-������Z@)]�Z�YpcB_�%�2J�U�_�,�O��Nh����g��G�o�\cly�{��F���Kg[����2I>�� �Vo��LM�P	m͟�J b?2���ĺ�|nd}1���W�e�=�����«��M|���f�y�3G�Z���~YQm%�OM8Ye=����������	:��b�A<eK�e ���H�{�c�GR���lƑ:�D�7�;E�����8Bj�!�B�sU���X�:�d!�iY���Qj;W_꽔���0�nƹ�.�6��Y�cCK�N������^����@c�{ϟ�X�Ԩ*m=���F�G�i��	�l^��I��o +�� �u�#g�=m� e��s��L<ZA¯<����,�^T��Rt>H߃}�ƅ��4�H�SY�{�3���:䖼a�(m:��+Mٌ�2S/Ԯ;��r�E�����+�[��l���.��U"'B5��v��I��5C�5��{��d��syXhQ��6����YW����V�Z�d2�� �-�l呑"����G+	4�=��SpJ��Ĩ]`��TJ ������ ��/.�{&���Ȝ��"��)�Rз0LZ�~�����Qz��t�ӠQ�Id��G2���iT���n^`Mfar���ؖ�2������&X�=�W]Ng~�:T��ͼ:q:��ZX�I�������}��*G�"�4�g<��Y���J����Eo^��V����Z��=༌ΰ�e��Eʺ'�/��a��xԊyN`
3�����E;m�k��9_���7�����k�I�?�!�^=��E�piHTml��
������?��/�tp?��'�d{g �n|���5P��eq��Ȟ���
���W��O�''2K�HB^����tn(�ޡ�Ef��|��>�1�/旯)}��(Xא���D�5��7��M�l!��tRt�'�,�W��R��o�nt�!��"%L+��v���d��p�.���p�G��$CM��D��u��0��[6
�)��i��#f�Y�S���B�bV�|\j�_�z�:����n3�*����Կ)y۷���c
�����^�$��t�Q�@���g��I��h�QA�8�(�Ƌ�&�Tk�}��C�v*�4+��5QS�mG�u�

.��L�J!�?-M"o_3C( `g�x���fJdD��A���+�,O����� k�6�I���B���E�s֛����h�>��!�OLXn� ��5up�8�8�wʡ�Ioܲהa�bW�qL�j�o0Yl|�+k��)Q��h��L����ķm�$���U�^tm��W�r��U��A�F,�`@�Z|�M�� �����<�o�Vge��Ʋ����t��9މ�#�	5�GI��L��"�*i�F����� ��.���/�n��E1�p���l�+1ٻ��9�d�58�N���>S�u�]D͒�/	a�Fϙ֧��JK��#p�]@�hӂ�zbH���Y+
������ �o���DYk˾�m�7���w}/��|�����	���!y����KU�N|�<���T�2��5Eb�?eOP�j�I[�����W�+LU�6�u)�:L% �M��%c��k�Gg��/2���	�Qs�ne��dť���r2��M�0u�:#�8�m�N)��ٰ��pq�l4u ��
7�!���xCb�y�6���˕�&$Z�u
RC$�`���Dc�o��`��p��,Q�Yk�v�����~$?�|��[�A�Y��|Y�|H%!�~�I����;T�C������&y�'���Xb��b�OP��>���Τ:qH�w�#\fB�PE�@�
;z[r����{u�oR�b�Br/ƺ�Z�#����-�d���-��/Evp���^��Ǧ��,	�n�֔ݝOrJ���A2~"/���Fm���ъ`+�=�)Y��	�'6����d��<tނ����� 0�O	�A?�����-�͚�����+��K��[�mQ���l���t������gP��y>д������@4��
{o��c۶+X�	]��{��U���
6�? 3��1�j��c��eA.�����#2��S����	ã ~������yX:<4
膺��q��D&��pG�z�����Y�(��kOV�.|<p
o�uX_)�x��9�@ס"�
�+J��o�f��|r=b�ijm�Y�I��s�|c�-ff�����6O8��69Qd�(*7���j�J�l��g��І�,�d�ŗoǙ�Us�[��]d�+�s�H�?���xs�F��0�?nXAEP�7Q@��=C>��E�S{L��}��m�ڳ�\=��{\��^,S%�B�n]��GG%�jQs�-�t������`F-�������P/��G�y��J������Ǿ$k�Ɛ����W蚱ً3'���3ԑtվA����x�C�����0a�~xe+y6�O {��4�t�?]�*��8D���(!���*�O�6r������E�px�����1(��%��z��W� ��-��	�4�/�j��A|V��6g.p
c�.��`��N`��f���)V�+7KvʊC�xK�:KT�I7�)��W�*{v@w��A�#���M[� x\.�ʳ�&;���4���e�ag��aEG^�{R��X���;ƬDe�xtk�Q��
:�U�~�#�?*CL�������
2.kЗe����r�*��y���!�`��i��&�c'ͅ�^�F��IYz����+�C���%�/0�����5b����CJE��!X���'H m��0�~f�,2��v�d�y��!Ъ��ćʶ��Q���@`Y����8&P��Y��i��D�Is_4��:��a���m��W�.�8M Z��U��Ba��M�/e��	4 �Uu���hZ1�I?�/��P�7èm�����[�W�mT��3G�tdqCG)����^!� ��)���F���O��=�v���'���G��n�-w�UI
�:\Ӹ(K��
� 0B�! �!%ۇ�Œs�1�������_��Ƽ�AM04xw ���莋�9f}�ap�7Q]�X^���f��ӊZ-q�R����4�z�����k�
�t���n�g{n>�Rݒ�d)� {I *]dTC�	`�®S82�dO�A�1��b�GA&@
SES��$nLv���;���]����};�GH\����f`��aT{�㼇����M�ŬK`��tB[��"�%��	R� ���<��������>��-D.m�ʹ6��{c-�?��PI���(�a z/gH�#��:��	q-�fe��J�<̌���C'�d�GlZV�kv�3��Q�q[*��j�}�V@����Z}IYA�W�^�Y�e��G����or�h�����>�;��ރ�r��ƛ�v,�Qxo#H�*`�aK���Q�2.Jc�ڃ������*��@���χ�3�����Ewݼw��<�<E�[�ݎ�sys�'.߸nS�|�`��r���1�[���\+\K=����I�C��f/�M�O6z�(�� ���s��n�g���e.�J�����W-o����3���v���Ȃ��L�^E��ӱ��_�]�*+��P;L8~����m9�O�s)�S���x�5�v�w}�>O�m��[���p��6`f���4	6}Fvm՞Ȃ�Vß�5���0?�]�+cnu��*�=�wSz�GD?G��Lzcl�Y�ۮvLa������T֑`q��t�R���,\A,�����]$������mDS�<��n\\=��w'A��%y��c#S�"������諁���#!>3�dRK�d�[b�+�x��&�N_���^���,8Sl�p_��wM��D�v^�b��D�Tu�ϗ���S]�s�4/c�ٳ�0�\�ԭdlC��Ц�8d������ö��Yrj]���oCL`��:|�C;/:���?���6�3��IWI�l�<܈���,�{�D��_3�M3A�/e���ހA��� @�[X�6c�=�M:�W�05�/Fy �x�����\� ^Z�n�1��?�J�T@���☦�Ě����mW��:�5Մܣ[����L[s/�5��e��[W�>��#����~C�t2C+;d�-��j}��fy\F�*���s�d��+@��|	��~Rܡ�5�jA}���)�!�%w�c�E[X��d=�.ɭ�Mj&ZY,mٵ�����l�rE���hb���L�N��a�q��n�
�s���*�Yݩ�c���j����� M�Z��w��#fF�<ܐ���\{G^�s��n�Q��<�Ջ�������|�����ꧧ,:��`A�\<�Q.Q�V@A᫇�ҋg0- P�z�G.=T�6�!�s�g�y�2;;c��,J���N�XlxV64EB    fa00    2640�7T���f3r2՗��<h��ORUY(	f�A٪�g�P�:�d��A�g��0=pX�Օ$1����rUG��:a~�8Nkv����U�g搓]��U(�`O��O���f�fqh��)އ��R��s~�iŠ��_2g��-����~�*�f�����k���]K��	Ę�C�x�ƥ�qn��#���r,��(���PX)�?��I�g���d�-2%�E+�$A�u(�����5�b�����2*�M��<]�B�f?E�.�y�?Yc�5Ɖ��̰��-o��.��֔�e<3�v)��$�ـ�5��Ny��p9<�֜2?����B���eqd�M���o�@��Co�JKl a��b"BJ�C{����m(,"��*�Nq��/��P�	}1r p�,�eSI����W�T/s3� h�����*�����ᕝ��o�yB~a�9Ɖ�}o�&׈6��Dc�o��xCۮ���ߺ���l`�af@)�U�h9�������3S���;t淺=��U��Ĥ�"�� ��d��4"`��W8d{�zvW;=餯l�H�{��8�,i��3E�ɬ@κ�fXN� ��"z�u�+�:5�	�dO�G�m\�3��v������������8��]��n#��^O.z&.W	N�j6�xlzTEk�s)T@����Ev͋wԪ�Fb_�B��'� ��u��w��4��q���k�4�i��hQ�Pw]<�`�uC\�<���'��a}e�	���j��b4_�a�x0�T�Sg��?��c�9��k^��j	���+HBfT��'h������s��6��``V��F�U@�e�	�l8��B�h�s�cpr�k(<LV�i{\��ɉ,{4PJv���s��G�O[m���Ɖd#�8|��+����d)-f�[^{�lIao�`F��i�Rr
�l�n�5C���z�j<!��j�dl��.�?h9�DQ� )���/@L���,0�M��1+�#�KY �xp/��&*�敬}�f�7N�����>�r��w6;ƻ���X��wP�8ө8`�2��y���>�A�M�����*y�ނ���@��4x�ʃ��b�àZ�y+!�r���]!�iSa�l���Jg�jE���Q�YV?g8x���Փ�v�+8{'edA�GsE���\[.:�\ӹ��YC�</$��P!w�$��г�P�����Î�����>��e�d{U�k���i>�̖'�짓�ô���W-����w������h�UKDl�IR��ʐ��jғ��8�.%��Va��'��ˠ7b@��~̽�O��d�(�R���u>���LI���H�-`NY׏f�G�W2b�6�0�"p;�^�Z	�	���w5���Ƹ��9PLL=�VQ:�T�a��`&�$�h#����kx>��#�6�"�<���vW����д�a|������4��{
g�{�����WMA�F�VzW�����`�9���Ѱ��0�1� �U��|��	:B&��w ����y�S�H5Cj���b`�]�,d`�4�D���J_0``x�al���?g�<�>6	PK���oT~d?��$�1��^�2]_�Q}�esC�� ���"�^/���Y$�� e�F9�!��Li�vS򏹚�	} ]k��������^�;���?w�iAqy狽�`ڳ��y�A ��(�p'K�<�t�(�[Hw������^ل�BU1I����2R����,��6V����zxmdO�Z�/��4���j������0c����!}�M^�o5:c�1G�ތ�*|�O��@t�������F��'���K:?���IeB]T��V�_�:�"���n���WhߞbϕuG2�0SR; ���ql���yt�������d�A9���L���	L��rB��nL�o����b��?E�iH�"D�����X,\�pdw�g�b��z�9lͻ�l��(X<�s�0���џ����]��̷O�=�Ζ���0i1C�ꊼF� f��lA���``�����2�A���?���?���Ɣ)�z]�`��'��X{������Y[Ҡa|�7B9�A�"�=���}ux�S�����,Y�Us���ِ�"+k����8���p�W﷦S`8kz0n�	?�S�����'��w[��_�F�O�[�S��;g���A3��Ւ��z�sl�.U��$�PK�����l������!N圧Ov��vl��=:$0p�%����辭���%��A��p�6�)ٷα���:��?���"�LqC
������$�lK�����^jV����uB�;Y�Z�
E�
j��*��B(:b��c�[�8�D(	���	O��?�����s�����[j9��[��!>R�ݺi�J�%����͑��l��o�r
��uES��m�ʳk<}�,��:{E��@-���������]���j�`H�Zjuͤ����<�:��~�������RP:���A/�����b������:e�AY9_�T�a���&@l���J{�i�dL���%q�Lh�)�� L�D��">������>�f�&{s-��y}�2����.dE�$_$��ű-�Z�ܙ���&���t=+i#~�%9��� ���Ά����EU6U;w�����фL�o��lZ��K��WcK��+�%J�ڿ��e�d�M�A��T�IE�=`ψ���j�Ϯ�ӣG-/����66�O��N�Nv�sQ���P�MߒzG��Ȑ>��s.]�)����x������$z޸���H�Ұy[I/�	�Dz�	-�C��gA�x9�-7����`يvR�$d�Uo�D���̆_�p��ǝ @���D�X7�
}P��EK�nCf�C�B'#ԉ3v�}�J̏;�����m�B�!�0�g�5k�5��C\�Ɏ1�è_����[�/��C2�4����׾�Y:
�3�����Y�ni��0�tRd؄��3PB�'�L�wy�\�����њ���i�o�W,}f�)'Pfz?FIV�����"i�X��'$����1��<3��>���?�%��zr��E�u��j��k�.�">c��C�8<;jߜ� 휴��5^�}�n��e&�o�0-$+/tt���5����0�I���+$@�}�������@W_��p�Z^�Ѡ���U)'|�EnWȣ.��8�P��S�}mƋ�ϐ�Z���	�� ܙ�=�,K̍R3=�74Ra)��,-�����㕒���2�k*��}�
c]�۞���V��;K:!Ք�B�'�E;���=]E���eo�b��pH徼�Yp���й�;�!<@y���B�L'G�S��{A,�W��Z�)i��g�>x(�H�,�@����e7�O]٩�����G��,��Ÿ��5�}�Ԩ���'�1��; ^v�00&3'��f;�+%���A�ڦ��Z�@-�(q�Xs�Ğ� kH,x�O���4��@,�k��v�R=cs!#P}G�Nc�/%o�6B[��7���2x
���$�Cp��r���0Cp�E��ǿU��Y9t�T��g-:`�:��ji\	�L�~�A$�����9�Ur�܎������f̟_`��M����j�GO�j�����$��&B��Ԟ��f'�K����ᨮ��ֱ5:�e�:�q��(p�e\$� ��d�\�۸�ū�|��4�ɔ~�S��TY#ʹK���vT����e���	S)�r$������)�Re6��"����>2<�ji�MTe:�Ę��9����p�vh������ ��S�V�4F$��q��6;s6%vފ%���z�Ĺ+Y��k'e�!I��>ٚ�W�*I0��A�j��D	���f#�d�>#�X�2�5H�I�=SVG��{�y��2�����H�3!<<}z���>�Mgq$�
�����=�U��jHb���?V��E������=�O��}da	8 =���.�T�H��e��r��[�u��.>�ɯDzA����T<�1��BD���cPO��N���ssX�;��#��ba�\Ax�#]�sė�]�u����y�<����N�b=S�+ ���P��Q|��7t�i��؏��>he����&����?:F	�:&�1?��ˆG��"?��U�_�5 `�����W.d�.��H��o-��g͐��V�}y�����E��ٙN����
���Q��&C��T���<��&�([_op���2}����
��9Vxp~'�7Ax��G���l�Y�8�V<L�}@�!�4"� ����i�N�n/���-dwש�������^���w��q��G@�o����Oӹ�Ó����H��~dڭ���O����*dgb�H��9�@Թ8��N����������4���6��--Z�zb`f�|Ӧ�!�LK�$���#i�=� ��	�
����<���Y}�.��ʼ��s��U��«�@��#���T�������S�	��?ۂyt#��Ϲ	V��V ?�By���Ee#Q�Bcx" �v�9��+U�q�\-fU�ĕ���9F+
X��ɒ^}5H&�J�2�`�h4�����յz�8�Px�r�!�ST�j:ȴ��GA󢀕��׊<[}�۰��7�����z�7�♊�V�Z3���,E`��-��xRL�=�w$�6���a7���}���w�tU��y��3[&08��]�Z�,EJ��T㨊����2w��˳$7���R�<���g~��d~8����W�If��ޑ�}��d:�Kp�*�>d�9��Cp5�/�R�L�˽鰴�0͢���.��@��FhW>(�*##��W%�X�wLj��s��v���g0`��_�h�֛b�m�$� [�f#�ͥUc����~R�� "�u=���s>A8�����Js��I�:J/�TLً��C>�2&��g��i�_�{��5]#i��X($E}Jr�:�K�D�8�l �D�����@��i��A^�IC�@���ٖ�`tk�Ƽ���hO�RI]F'moOS����s����y�L�4�hsO��b�݃Y�:cs�=	��|�Ky�TƇc�a�A�+�xB���J{1D�mW��lk�m�ВC��� �L	��0������w��?qp� ҙ�9I�,͝�0��iR��:���4C�qIt�����>\5> �~jy���i��쳘#����`jNY��,-�)TC#���**!��,x�Ԁ8	�Jɫ�pg�����{�MYk!��2�zη����5��bV��b&���� M/l]��^�CΨD��|��xZ���y(dL�����i�vlKɒ�EI#d�j�L�`bH��K0���0��0���քg+_�]��h��k31R^��*��V�6D������ŞFM��C),����N}	c�'����ʩx@��F5�_i�����8�à��<�����RQ�:�S yn�+�wu�t�6�hwK�`�:&n��Տ&x���f̪���"�k7�sdWX�Xr�<�ƾ6>�����L�����b|�h��x@+�����i?�Ϥ���gu�]��QQ`k�,�.td�/X3=��(>Rd&��%�2�>9t���Lr�6��MͥT�s��P`vƵ�c�Τ��lji8Rs�(Jv�G�M4�b�cY��7K¹FF�o��x,��7JTνq��Q.X�X;>Keؓ%�|�eF��h��<M3���r���������7���^�7"]UY������m����#��r<ē֖����s��S�E/��������Y�1W�q�콳�X���E��E	v���X�D�ߟ6��s�c,���v���JNt�@�uO@���P�@��\��7����q������6k��!%����h�/61m�e�S��T���.�P�k���βq���f~c0���� ��t6����S��p4�8A!Ӓ��Rx����B�V��0#M7T�ɋ�թ�������RH��n8_x�қm�d�ߞ�ᥳ�{�o?�܏��:��@z�҂��%?�:ø���sϰ������Ei4j�5��~%q'{_ot��f�>s��W���j?R��ގ�S��%��̌��	��j����<,�7����.����/��]�M���* ����@���U���[L���m���To=�����X7?`�0z���#�_�(��$\+�E�Ԃ4��*�޴���4Z{S.�+:�� |��|W!����4'ˬe�y#΋����/I�3y;hLd^@��r�wG�#�<&�RQ�82���+l���8�-�!+e��8z��e2��뙐�o��R����joԑ}3w㩐�/9Y��)�E�x��d9���B���>|6���s��H��Rae��� h9��L����ZD�*�@>+i��#��J��T^�=d�J,�v~l	E������",��e�rD�ym�bl�ʸ8ˮ�E��rX	��P�?hn-[����}ж0a-4[���7iE�m��e�3���8=�Nc�8P F�SFW�I2t?��}��ҷ�UOB��[�xP�?�%���(<v=3�25"�0�]��6�DXhp#��U��4ݒ[]�'nĐ6�V�ݧ��+�M��茞�1!CR�CDԅQdE"���y����:`�[������_Ƈ�B8]n��5"�{H�y� ���)�Qӿ���IB�,��vu;N`O�)غ
�
��)�����Ǽ�e��d��4��@�7o%�u�Pr��"�׷�.��t��"�i�+;�;�ߤ��I�pQ�5F���ŷ�_yP &\֟ vq顆c=:n��!��?'��k����8�R��lϹy@�J!#3|v5EP��D�&��r\��ǼU!�ߔ� q�&���HdRٶ���KU~K*��x�|�k@k�����8�-���i��O�ua`ߴ�}JA�_��24d׽�a�NGV��8��d2�ѝR���w�Mo�.	�`�����d�Jc���L��uA�g�c��9̇G����piBWHڅ�'/!�/4���~~�|�)AD�^�������xP��`��z�͊��#W�1hU������ESoSk�|�L�P(j �]u�(��%/�04�Nm+�v�/j-����mQ&R�dU��ă�e�����?�������S�2ǁ��'9�nJ/�nuB��.�2Y�W�X���>t��z:\��������[-�c0�B���U��b�O��'�����ʉ�\Im��f)���q*��,g"� ��1�<�=�|���{{�Ҳ7+C��<�d�L�+�>�-��:X�i^��P� ן�"���ţ�[$����z��1�v�<�&)�[��[���ٝK�Ȅ���r�t�=L<�v{d���X*l����tޢ��1��B/%�x@fm袜bF�JӲ��D���q�ʏ�jS�hnCcL������Jq�>�����c��@��]���D7Xi`^zǹ���$%��!�D����л�.����w�����n�I;�ꑓ�{'���9b�Pv����t�J��8{(ë�q�<���8�S�#I�% ��DpaRj�b��vx�\�#t�X�SS2�eHtq*�l8��x "���?@B��\�= �f�󙆋d�iB(����lg.�c7y���%�y���ϵ���Sc��z~ X$��k�p�k���0���j��;4�R�*�����ͶxF	d*`���#^�UrL�S��]hn*�Ϯo�Ƭ�=|Ԓ:kp(8�i݄���ou�n���1AQ8��r*C4��]��Z`�G`���~�xJA����y�ۖ�o�s�o��K§������~)G=L�|��pM���I����Vź�\> ���m��sj�<���@�;�">f�8������l�"W\X��@��O�qc�>ٌ��� �&/�(~?���D��hHp�H�ed���?h��o�F����+�SX�'��fc� ��+}$�W�o	r��-�����c�!x�
��.}���u��5x��X�|��&�_V&"ȥ��Iy7��Z��P�k��ʾ��=���w�,��L��*5�䟀��(�o��:�9B�ύ�2�<��ę��K����;ʴ@�̵�����y��=it��ȯv�V�F
��`�]B�Ax�^M=�ޡ�=�f�@f��X&Cq�t��m'�{�<`��c�OR򤱟��XqI��c��R�r7{L<�6�G��M-�9"ĥ'����po��\h�Ƒ���P��1�嗅Z���`H6�OIA䝈4����#;���/Ja��R׬=��o�K�q	����ʚ%��
F�"� q=q|ъ�O�L�\�zB<E�f��]��Oi�LAք���<�(�/�@'H���9EG�%�qJ�{�A2	 ���#�H)vB�ք��C�k{ �����]��=�$��'Y�Ҫ�peZߘ|�-T����6��a��B��` '�����\�Uݿ"�[�!�ŀ��&�X����6�#|<�mȹ*W�s��xfsq��󺞴�Y{I(��O�SI)���	WB�#&i*��97Ĳ�ƷsE���{�%�p��0M�oN�P!5��ή�Ik�����hnW~SI���w�!�Sϒ⬴I��o��|_�C�Lt-eD�:�j��"��{��͆*���/,bB�����Ž�8��rq����a�{l��U&�~��(��_"p?��.�e!�,�oN3=Q�N��.�b��HZ6e��4����jW�5n��� �u��,N���R��[����*շ�
1�=��&��%o!�;ZzRc�k���{��=�t��c�y}GY��(����>�0��������	DD��3hJ��r��X�<�"�QϦ
 M�}��>9-p:`
ֶI.�H;�Ww��o�\՚�d��;�R�'?��!jwr��P̺A\�N�Q����%ܝ���_���:�� �0�H�A�*�$b8��}>��w��3u���[�.<hX�.���5�.`L��
vD�G#���ڧ�PY����W1\d��b��i�S��~���5�����l���N�s��J����W�����7�:��u2N���1f<j�Q֘��4� }o�����7j�DC����I��:��'�#3Ud�'1��pe��Pޏ����EP k�-����0�Y#��b^�s��'���eL���zW�",��yP>�@v��ɴ+u�D�v5@����gw�X��m'�z[��w�Ʃ����6Dfd�&�&k6�5��נÙ\A;���[6r��GA���(1��E�s�µ���؟��6D�[�G$�9�J��s�鬒��d��F��5����uꩵy��x�M$�`�]�Tp`�e��5�џ��q��躳_��3��!`��gkS��U�e��]���{�4�9���+.HQ�_ش	'gT�=:�[0@� �4��S:5 �6	i��S(:�rǠ�S�� �r�N!�扖��� �J��ڠ}��fo�y��Ɗx��Yã�he�Ԏ(�9}`�Ų�&]�M�nC���!M0(���fx�]�-d��j1���*+��S�i��*�E�1���"��E�4�/��;�@��Q�B�;�>����ƃ���2#:FQ�:�&j�����mK��}�<,�zZ�Jm"�����0�����L�q�peݑH��"��XlxV64EB    fa00    2680�߶x�B�TT���s��� <��8O�����C���e��7�`w�	>8?��f�arE���yA1��W���F�d����MUf�Ÿ��x;�=3�v"����jw��5�� �s9B�0�Nz)Ð��9���+f*N;Țx�u����i��rŁ���fbt�H�����?9χ�RU0)&7`�IM��?XR`�i�Ej������������CXeЃz��wR��هϴ�m�A��L0��*`�x�/���Gʯ�X@�h+�>FU1q3�v�I�.e��{�Aq��X�䬔�5���	ڗ8ċ�4zop7�Л���Ew}cY�A���K]���Ҏ���p�
6�|��^ʢfQo��{�g��,��w)�4��IA���I!�$䌢 OVt��U�(��n���?i�Z�^�Q�a�an �̱,��~ZxmLfѥ�]����7��X*.bB�yJj$��S�8�Bu 7��D`���Ig:xΪ����v��vwQ�D��X��ǌ��s*j��¹=P��Dpg��su���Z9��QY��!ؕ鮡g�����(�C6�Q���i�7�X�+��1�$����@%m�-O�
����Ȣ�I�o�8���Z� ��y+�?�\�啬�$�Z=̕��:���:�x���,GO�G��w$b����:��CY(�G<���J����F��G��� �?q�W�o0�ua�|}�<�:&R��e�����HT�	>p P����#�jB#B$PP���K ��z��1�o��˫��VP���c�B�36S�B-�z��bC^����aΏ�E�к��9�fJQtA����}���#o�)XzTG�'Z����vo�$%��4 ���6��mM�`�m��An��G�n'����j��eXG���R�^d��2���peG�|oF�L�V�����,m��3��K�h��N"��p��'�{�FdwΕ����rU�̖��H�+G�Q��S�(����͋��[�2v�ӛ�&u��o�
�8yq=�7R�={���T�_ly\`-- �*ʼ8��s�37��(ˑ�Ń��+q��v��$���,����C~�Vr'�뱘�%`[�q;K�ͼr%f����=�c��Z�!���3���8 ՇqF͙��ߤ{c����01n��v�N�,}��E���!�T�t��dyAh����������6�����h_9UUY���eD�1��)��o�V�G<�������R�^q�Cq�6�%���na�*g#ʂ��]p�Z���e�<�p�"�0�OBJl7��q�FQ��R��a� ?�6��C�J� h��F�)K&��ǋ��~;��*!�)��,�޲�
9��|�ՄsQ�4��"����Tī�|`G-�߲��ƌ��m��aiR
05�$��s�����{�z_!4��IB�WHޟRZɑ�;����$�J_�E{EX���6G�ea��Z�'�y/Q�ORNU�#��Cv|xJV���,�Ã��/��)����8�GF�kP�KW��I�N��N���`�M+Q�K����ږ�*龺���h�/���	��dO�F���@�7��fmx0z{�H�Ҍ���!?��Ȗ/4H�$�0I�wS
)G�ҁĀ�vc!�f���#�S/g�Y�`��U �d��܄o�\�1�UB�陃[�����_>/�;	4���[��1��%9���k{�q�T�ǜ��@�CQ��[�شm2\�8��Y��6�ՠ ��C+�.��1\�E(FJ�fRI�WJ�?yF�8����
҅��N�c�
�:3���Xʦ}�=2��c-��P����G%��)��ucKKXW-~ �zj  S;Ӈ�~JC/����9y������(�m�8Y�;?�y|��1���B��Q�B�9��,	
r�*g��~%�>���Ǭ\��."������X���c�f-��Fc �_,���X�k`O|;�~@jDW���&y`���jO1��}���Sg�7Mj:'Ǵp�����9��Ԛ��@@���"����؏���;Aeg%a���0�S�s	�v��,;(L�v�#2�W���Y��FΉ6	I��Ivf�{X]�W���|�/��T�n4��Y*F�=U�r�I-
R�W�cF�*���#���h�[;�:���D�S����R(S��)+͞I{�X�^�O�wq�ĿDj��i5~�^Wȿ:R�k���E&J�XAInv�=ŵ����	�T�Y�è2Y�ߗ(�tH�����k��Y(��(�bYR�}�����4��Yr�Tqǘ� ;��5��p*�]�������s����2�3a����is������Ɲ�G?���5?=����yh�F����=�)�7V<�)�1�[P헭�J%�m��������D��ġё�O�!%���@���_�Wbi��Pnt���3Ҳ1K�����m�/#iz�K�x ��'Y�c����sv"���Ѭ��ݝgy��t$��>��0���,Y%y�H��m��3P��nV8��T6�)��mx�x:y�	[y�������a��#��Ϧ�H��D��7-�Hp���'
ʢ]Ϩ��e��B�K�>�jBDfu*-�%�N����r~�R��cD=-�*�է,�Q`�6��6���ђ���vI�5l��W��(�@��j!�ؚ[[�u�yCs��*�D_�~�s�[���e}7�� [��Y
_ux�h8e�Ց�}k�5������`��c���!�*�5�y�10��8�B�C��
�Ulowa��ucsB�ϕ��Z��=sPG�E��ksp���A��s\����`/XǡNO�����X��#yʶ�T�fr������{�L�P�P�(�|�wz��"����H�ﱖ	#1��=��d(�V�5���(�=u��\�,�rC
�\��<q���=��J��@��Bó��4C�5�l��#��8�q*���u'z�3U�6�[�3���^�H�$�.ueCK���ޒ��Ry�ޡ�� D�8&���a�<��7��'5qǞϲ�F���q$#�q�ۑ{d�1�	������3��A��� k��` +��=��oM���:�-;< �@t��	�B��?pn��7_"۠ʱqH�Iق�A��kp;�2�6�a�Y��{K�c��0�:v�b?�x�ʃ=w��/H��U�$6 T"�&�[���M��彞c����*�����|��]2\������.����"�;D� 
�������G��ت@ۿ�E�6k2�/��o+^-#��{b8g��I��q���b�J����8�^H?0�m��r�6'Ƃ��v�g=Sx%�ycbe�E�Q��HFp&K���J'���dU[��}U6% DbY�E�ӅЀ�c@��X�=v��!o��R�L�|�%1�龅jƵ?B|�Ѳ�9oJ�T�R��&��u-�"���#T�o�����8�*$��Cϝ{"�;��{��lǙ�R���#f=�^`ڗ_}���2׏�3�P��b��x?���k�;o�[���w��^K�L��yV:�d�R"..Y��"I#�MC:}���5�f�\	�J��O���+�L��=K�i��KK��ƌ�_q+��e�͚Sp��éd1�P�M^ˈO�N��,�k-.;Q�9h��.&J�ml�@�3�jdf�G^K�sV ��}{�F�&8�7"���5����}�d�zL�)� ��y]$Ŗ�u����/�[R��9����?c�3�����d	����/�`��[i��V�3a���i�O,H���h�G�<��Y��̸7�3���D,Fqh�G�`�q��Q02��~�R�{�����̤�q�/Z�f�]�N���b��"�ʛ�v�Db-��P71�X2D��N�B��*{����0qƽ��i�WMkI���Z5ll�?�+��ǈ�1�$����2�J�|FZ�8'�؏K3lR>jux��җ�5/OV�D^�n���c|O�$�MՍ�oˢ2"瀀^��|		=�
H�#h4���Hr0�&�3�~�B����T+���5|��x�����.��]�!��k�593�8CA�&����B5�8���.��ܑ�p�C�̞�����!2��!��U;j���o�/���k�����*������h���"/���� ���Tow�ұ��u�|�m<(X-&���ӄ?&��1���]ģ�W6��ծ.o��ܯ0�l�;ɅX�B�|�Yr��R�����=A5ZiS U�zV�b8 mw�/�%�/�{��-=M��6��F�$� �	s���;D�����B8Qz%�_۲��=���w�\_����Y�w�5.�\|�础�K \|R�+@�Mp��@j&�P
�A2�W�4�8ϫ�[r�@��[��XO7ޜԈ�)A��o��Q��L���o3[����_I�5��wއ�&k�)�8L ��T/�H�퍽R�g��5��Y�{�Q�bf-=�%+�.�g	�5�Sź�W!5�a��ă�qL<�,ݽoO�*<c~�PM͓X�T��l_>�Lޮ7ԕ���Cx!w��׿�M�ߌ�X�\��<�AϤj�V���4�(�Dnb�Y0��Z��=�?�(�Q�
z�=�Ҵ�9��*���_G���㤛˶v{�U��z�&Io�c���&�´p3����k�G�V#��k^J䚒�t|��G�5����mRռ���o�p�2;1a�%��
�p�Dt2�$i�����Q	�l}h�ɵ���zS��բ��c?3��(t'�\�L�r~{<���O��c��/G���svqr��>|��|7(��`��k�A���]�<�w��^�5SB8Z�8����銤/)�}���w0rP���Y"p�M��ϙk��b����2#��Q��Pc�q+������<��*AFVAc8�$w��,�������Y�H��ώb�~�)D;c'Ua>x짲�A�c�x�m��9Dv�CMC��;�VK�Mu����@-XF�Y���*�^ۯ�L�SS�Fh8�VLC|���:�qu���|��c�,48�<[�R�]��khz���h���p�xn-{��O*4
�8��ޓ��2�Z m}����poV\D�I���8(7L���q�W�b>޵NR����׿9 a��1�}Yҍ��^m�Q�ټ;�t�^[3�n��Oi
ʍE��d)�9r��n�*D�7F�64/<�&�W��u�9� G5����捳��+��F�]P�o�׆�}im��ߚ�?%q���M�~���}�[��Cx�"s����?R�ݑ��/C����ak����J	�5#�t=%��՘RV��+��J����}0���S״sd��LӜ�&kd�k�r�B�E딖��}K�	�u�!�/eq�? a�P-*�@�&��#L�ne����J#��Թou�o�
J��,�p�T�AU�/.k^��SM����]�%�����h4b�ӵ>T�0��f��Cc�"�u��n��=h�Ҩ �H�b�) W�Ų��-�o��-�?�����P1~�ڳDg�����U��MWx+X�Z�t%�}Ǽ�>�x�)�\|�����'����=[~��E7�����&%�{A���c<n�x�\Oɲ�QeW�`b]�>I�Ѵ�w��Žy��#1�a|z�:Tz؁}���K{��7�;%�����QLZ�G:��7���Ό�*Җ����rjov�k�w��@ㆈ6�,�k��t&�k��aR�1��u���2�]'�r� isէ�C�����EP�0H�����/+d*s	T*�t.�{v���\~k�v:[�R 
B-��O9����ؿ���B����7Y'%���QK��A?���CS�B6��I*h��	
s6��x������@a�{o� P�����&���E�#hj�|��$�CA�G،��pF������5��+���z��~����~�]y���!M�EJ%\6�dwW�r&Bג��D��҅�9�RU��	���\8�d'I�'.���C%��Ϯz̈́@U}Yvc�}�k�4��������<��­G+�M:Mf"	 ��j���-%a'�~�졺�������f�ن.J�m@�w�8�ixQ��e�@9�����' ��e�2Aa�hǳ3=�d��Q��˽�#�ܯ$ �V�CI�׆u����t&צ71��S��Z�V:�F�|/f�xD�d^�=�����s�1f
�ijЩ�b,�30.L.���_����:r$��� ;4��q��+H���)�ֲΎK��������Dqؕ�L��H�uK5B��J���� ��M����b�k.��	d@�&1&�6n{����Jg~�J\<�v�so
}¿���]v��rL������ǲZ����׮�l���~���@�Nw���}{
Kq^��G3�y��f  ��I����t!0�т���ya4\=JL������-ZA �6��(�sq?j�P����.���/�~v
�� Z��|z���_>�:�2y�wz�#=]"m_��s���!�#WV�-��r���҄vRyG�y��Ef��+jt��G�l0Ԉ�����`��pP�h�a�|q�B���[:��%�ӕ;�45���|�qۓ���[�S��x?�Mf�bhY[fX�vwH������Y�,B 7n��}ءr������yI	؎8riT�uZi�1�|V����p-������0J`�������Cf�+�Լ	�$�ڰE$/PlY��8�ukY�L��u�=���t���| w��r�l5���W�MΪU�����v�R� �d��Qu�j�
Ԓ�R��fa!Y�B�nP�Y߮^PwUA�U�Ձ��^ށ��W6��f6#C�@���*鲟�
�=,��0* ZW6`����:��jv�Ck��SGħ��
A�!���Ԕ�@M��Y�=ͷ>8?;%�K ,'��P�X�,����
3����6������ϱA�wT6V������Z���}������
�ӱ��G�.�׶�UuL�y���*l�e�Jؑ!ތN��`���)�/�-R�7�ft��7�b=E{[���Y)���T�o��U#�=|�  m-�	��nS��"����5E����� �WG�����z����b�O��#sa�"�s��Ƙt;�D������6�'�\�S�o(8WH9a�پ���K��9U)�GN��c���C9�+���흢���g�"'��-5��#_0�����\�Hc'H�s������\j� QL�^��
�Ԛ�OQ�.�K0�WPI�M~�px��[R7{��ȟ?3"q�m�x J�c��cG��Sl(BE��!�u �#yt��ߚ�S�EZ�=�k?z�@�$�-�̷k4OS�-�A�C
����!�!$�9V�@�:¦,X���^q�����=`mkb��N�AF�ۨ�h�`_�U&��Š�����H�RK�i���63'_�.a4Z�OW����`��Qꩈ�ߩ�����̠�����������cl�f���U�&w]M0��O�y�O�2!6S�:7O�>���.J.��p��ͫ���L��z�z��c��;q��N@���{z}�zWy��Z��vz8�e�TVm�N�`ak|7��I��Odf1:��/X<���X]�$��� �n�NqC23ŧY�hR��3�]���l^l�����{\���={]�H�M3�ު�zЙ���H�V�9I�.o���f�h������Y����Ǵj|#�q���,_5�D۔Q	L�PTl Jy~��z^��4]�?wVt������OP�e�Ys���AnL���+���30Whf. ��[������H7�\�},�zE�ڼߞ(�(���FߺY����k���+V3
��nPd��?�(��1�.�U6��\���G��!���[qR��-ʩƒK��^��h���f�5V�[��?��F��*���P
=�/�u�7U�?;.�x���w]�����i���ג'�&�����#hh4\�荺#�	�}�f^a�]F�X�R���\S�O��S�?-x� ���ёa���o���+���g>j��	fGw>�VN�zǡ��B]���+�8�������ɇ�:K\eg�����0�h_mK�-�<!Sg��˕�r|�*��Q�,~>��6���(N�����A��lZ��q�)`�!�-����T�?�� �3n�~���d�/Y�+�!�M�P��K6ƞz&�-�T0��Qھ�A����FY���Q�"�M��^=s���
�6@YG�l� �b�6.�d݀
��}��C!�r�!�w����L�9Xő%2?��*`\�)��P��sG��pP��l�)�\��t���ν�{�Q���pӋO�(l�87Ѣ5;��l	��	�3������܅�����3���e_"�����q+m���i<�Dk�a�ؤZ��>�w0�(a�/-��_�׸F��c���[�Kr�'D�F^]+AJC��P_���˘NP�,�ߧ�n�b��~&����Dv����y@���@�;��7��o������F�50&ŭ�

�����6��%ӫ���{��E��V���K�d0פY�7;���-�m�ۧ��%�����e�M��Z~�k�77�k�d����b�'�ɪ�f���F��2��k��6���ZT�<g2�Rk�ta3� ;0_R�w�j�/~6*,�z��X� �:���r"7����[P)�eP`/i��<��x�yp���P�up1�.�gt���rt�9��#���:E�k�6N9G�R���$ߧ4�-�5�4������l�Q<���}�"��rQ�K�?ix�y|�C�I���]�Nl�c����q��F�ԟ���m�yk pŤ,��W��z��>o/rvy�ѹC��L����d�N�*[�D���"�-^}-�}q����`1����le#��N��J�|���)E5	�d8,���Q�W��t��0K�9�fET�=q�e���7�A�AH���f��#f
���-���P:Ed�������B���C�2S����&V��C&C&��ɴ�+� �(nKrS[��&Oʆz�M�ߐ$��Y�_������~�x�p�KbȪ�v�"�r?몲.�E��˙��d9SU2?K+�)��;�g	Y�d������k�>���y�Ʈb���w��r���.�������G��1Ӧ�!����(�E!��o�U�J�EJ�[�;�
�7����5���Z,n>m�N;�ϳnR��Y�A���4w�<=#�;QO�"�FP��V \����"t��O��:��e�U6�XS��n��.�ר�sQ
�}�3$���|�N����i�G�X���V���Ie���
!�Qr*1����BV^-s������`a����Yno�P^��M[vR��,��H�nm�+GǪA�؉C��0�ORM���O&�"Ew������T2"җ�j�*��V�0ԾK��)�*p�>�"�;�]�D����:jp��Fy�+�K�ˏ��'�-���  ێV�������u�԰_�?ߺY�"0��gĨ�yW{�Fts�=�&c�KOsʵ�I�O�����=��>\։g��Ӭ�g�ugƻ��z���X5�w��#	�@��Ъ�������	����kM|9$�@��Œ0��o�rX'�)3�4X�Vq��n��X��X2^6�5�X��k�_�:s���[��[���]ǐ%:��,�q�Ϯ�꽛.�b��XlxV64EB    fa00    26b0<8�7Fj̢���?��2����$[����^�z��_����G��G�',�{9�����Tt�g��֊d�X��D�|�Ռ��2����� "A^U�1��� ?9��x�N�D�v��Z�����Z�C�'񞒞�S�:=�o�D�d��ޙ�e��}�q�E܋��Cx$�{�� �����Ch�R�r"� ;iL�Ϗ�K�x�s%�z���˰����rp7�z9�g?T���[A�nC��V
�Hiע+�����	A���b��ĉ�}�J�LJ\��{�A���?:D����N�P7����bB�⁌Dw9�7��wxc�r^�تA \Oi����b�J
Z�0ȳ�����S�<�u�J��9K��:�}C�	 и"���/ ��!�t�{W�*����5:�mûd.�����*���p�G�_ᨩ4���PJ�->�K8(�.)�e�E�>�d]��uݟ,���r-=E�Sn&�scT!8���5p'4E���I��wh������߭�`�YA}'4+�NW� u@0�S���̀������$j����$|fX��E�n�ϡH��Y���p�iË��s�̝1�nݡ�t!����螋+�Q/�3�3})>�gI��olG�DA0@o�SR33�?��wk�C�����2��H'~���!��O��d�9������p��H"�4>���E�|#�ۣYDA�ĭD�M�)]������bɒ����o��{9;b����(�\)m��l���N�=�!��xqQ���S�'���5:L .�l���'�.ӏ����-z��bO�*!����������y�`���B��z���Gp��B��	T�Ѩ��5K
rv�`�a��։��JF?ƛt��⳺@�8��0W�˧�[%�C~N��nW�����*�ʀ�bc�����Aū�}Í�M�����i&���9�<�l�uQ�E��*��gU��"Q�8�k���`���ܯz?1�#�]WQ�s��b��ϱ��Z�n�Xè#��P��e@�{� �M�\�s(���>�����"���c53�(�8�y���4�Z��]�%���qh�~j�y��	#b�uh	f�j��"vV8u�Rƥ�+����'<�`��L䏼Ty�2�VDJ��_���=Ś�gW���=��͢�N`�5���ݒ��V),j��*�~fn�0��p���i)���P�i�d��h��O9�au)O��w�Ֆei`��|�`(i���k�}�9�B����o�-v��	�(",z>g�'pS��j�A+��<TckHF0X���sE0Dq�~��A�֐�(�q@��^Ӌ	c�ٹ��a�,?7��&)_3�N��r�44��*#���ŪA�-�9�&�3F�ipn����c�0�� ���S�Be�i
%߇�D����r86��2w7����&_ЉoEl����m�{�l�苅_&Fփ��Se㶇Aݬ���t����P��aiK24:���
�ɑ}�d.3��EҌ��D@_ú��޾�~w�Y�,B�����?�����jSB��:�
]��[�V���(\��#�d�L!�w�r56ra���l����3Z�we��ƀw�-�g�G��vK��s�6G�K�Y�e	�U}��P:�Ju��&�U)*�DAekZ<�����_����u����E��,ݘ�=�Xl�m`���I�oևnh�0�.e��b���IwpޜsO�7H��
��e��u(@ ޑ��2�Z���v�A9��J��ވ�� ƪ�6@�Z�b`\}#��?Yͯ|^��s�p�J!�.�V�鴖1^�{����G
��`�xWg�=c�K���+��H���"�@�
i�~+-���	I?z�L$m�#s���Bt���hZ%ú|\T� �|��@����N	�1D��o��UD&�?dJx^E]`K'�rICCz֍Pqy�*S"<+�K�U��!!|�@e�b3ϲ��8��6�ʥ�y�ށ��ge��@�u]e!%����2��m�<Pj���\U �H��8�����U�06��Ql5gܴ�$���Dɂ[P\���cD���B� Ǻ���3y��w�픉�DH��<>/tm�]X�م^g����ើ|���R���e�,����r�4�c�3�nJ��lU��iG)�����N@6�4�<�������K�sv��bd�k�t��Ĳ��:9��n.�-+�.�K��Xt�)O�IBQ��ʿ7x�Y�\`���b����Z&S�El~�E�KJ鯰� �
z���ʃ�ń�V��Z����S����D�[n�Ԙ�0� X}K��SD�/������G\��ۀQᢿe� ��y`�&5M�軇��d`�T��2T�T�H�������a��&���>Չ�#4��h��m�-Mp����q�U��j7�=�[�m�	g����AaZ	_Y����\��i�Ro��2�놲r�0LL���S�؊���w���fMh�� ��m���5����$�{N�����ӄ�sWP��͇ �8;��,4�`gg��F\G�p���J=��˖/�M���Nx��[�����3�1��	-�ZŁ�B������^n�%V���h��J�}�҈��A����o��\��PB<ZPw�G��
�r�Y5����ű���aq�S��Q��a#)���T�ד"f��)�8��~���R4m�c\2�F�������
�/�ʳ'T#l��h�hX�&vP?(-��O�^år�jK\�Ta�p`��j����B���٩�����4�d����$+J�.gH~����ܭN�9t�D�r �=�X=��	�څ~p1�bqB�WG���+�Jë��!�O���
)��Y��\�R�,��\S�͍r���X2;�`٬�@�ϔ_a��|`��0����Y:bnU�aS��d�зj����o��^�=�j�uP��{:���X��p����&f���pe����
��)p��PB
V��t7�S C��ժ��8,� �)d�����v��h�^�L��ͧ+Y��x���Y�љloY��3E���3���F��:�%*:��^�f�9�xW|�T�UU�ʻW�%��*�|)U�{u��R�(<��X6�ܫ�j�ć�3���v��|+'�;��5�js���Yqe"�//�a�O�����f&�0Dm�l���%L�ѧ)?����Q1
̒?k�� ���:f�����_諾R�b38�C�o���}��I���I�ҥ�j�p	�����z����T�D�x��H��S?��py��J�Gm�w8�kx���.3A�.���AR��ɳO��ct8�uV������Žc����N�o�9�b�_�_������d� ���!�=�����]��$�@Ҙ3Ҋ�s��Z��ϵG`ɑ�Ul�J�?�U�8�p�	O�-?v�U�D�$�k�{u��2�(S"-�?:u�fNp�Uw�Y�ر܏wT1��{3IRê��u�E�3����	<��D�^��3�E���V�a�r��#� �C��G�&�y���k�uF�n�'*n�yZ�I�Nm�$w�a,3�*N���+���i�s#Ά���*S�Ǘ/�o�95)�	�>U�!�H�ә��An	�|c�'�����`�o��4���YP�<e�S�GQ�a���Մ��2����ץ�fYF��Qq�-�]�3=�Y�㇦�!���%�9װ�����@Cֈ.�`ۂq����`ZHH}�l��OrV�i�6l�����趨��:hn�w���qS;<[��2���r��i��w�3�o��'|O��0/�&ɱ0.&�|d�-ip���!^�/ݻ���w�sڝͦ	8��&튋=S�#l�^g$-�殹��ta�d�����?ھ�pT�+��V���ȹ��=��3�W8��>>B&��)M��֏�YW��M�e֢�'k�[�z�uu+7�rrv�*Za"�kZE��>6���e�5X�Y�[���n�J���9^���w�ˠ��
mm[Rϝ@뷃��҉%�m�D���WYU�l�d�[�DZ �j�dl`0��>����f�*�k9:x�A��#}+���26��M���
q�]�5�Bkfx�ܮ�B�BR��?�>���X)�����Pc���A������N6�_*��~�CYv�h\<ρz�TK���F�w]�$d�>��&�u	Lс���18�]kBm���V�_�Z�.����W �E+[E w���ֆe3��m�H�g�:A���x�t�0����%����	�A��}���@k�Q�pK;k�Ӕ� kF~��s����5�2�QF)+	�-���t�}7.N A��%�uCMh���2ǝ�����6V�L`\ʆ�Uʼ�^��l��,�4n��H�x+ʱn;�8�����}T�Q*�#L%�K�����������%&�a��.�Q���R�wc�4��?���C��'~S�PY|m����h�[�����3���ϒ�j�g|L��5^��M_�V�sW#3-�s	C�\~}|��B6�	?%)�<��x)P�O��� �|8@3զ�2����c.-e�ݣ�������Ƃn�V�d�ث)����%�oI�n!��������?_]��1�vn��e�P��kπ�JUt�-(�o��P�;���}i�r��.կuo�WHfֽ[1�א�<i�����|�/����r�Iy�k��P2s_#�V�)ȉ�� )�X������b*�����)�'��,N@����5���E����0I��z�8�����N�����U���\Y���)^��)�:�1c.�/o�0|ټ��)Z��f3�p#W��<�<v4�΋���p���7��C���a�H�,�F����W��0Pbt��z��X��jD��x����h�f0pN����̔����u^.�H�����?��fdr AS��v��N=WK	�DG3��C�jd�]D�����!�P$7� ��fګ�lYqy��I\�Z�q��#�A�3�m\-JN�P�x��ſ)w���<&��u�c4|����a�/P9`��Ů����^;	\w)0" 	�A;Cpx�������/8`�,��f���������z4
<�(��ׄSk�Fs,�OH)R�d�R���ݿj.z��'�[)}�̚i���HE�}�^��� 0˶���+��� `)p� ?D���Y����_����3}n䊭�"��� �=+�h�T��Iג6��}�	�iڨS���z`ԁ��پ&�����ũ]��2C����?R�|����e�`̀\MM���*6��$��3�
�w+�o�\����]a�`W/����/Ũ��n�%q���:{_�~
�
��M`���f�R�xՕL����!�'B��,Z�d
�0J�Vh�˪��� ������C�g�*�6 l7?+�珫��[a��	��� g@w�6��_���v�o�w�ΰ�4����?�O�k�v9����=����:i꿬��4�2a_�3>2���,�����d��V0��h�_��.�VS)������B=�9cC�����d���}j��3�s�$��y@�Q�R����	V�����@���]RFU��ӵ\���Rݤp�Z8�����O`�a[MqTXdꌚ��ϐ$�kp榚x���bz*���A��V�C�=���2&ڬ��T�+���%��]���Ǭ�Ў�
Htrz�C��A��V��Q����� �J�MוG�����u�{!��ˡq��B<�e�ww:��<��G��-я����S���tS�~CF������	�G�̞&%� �Te���r4��7�p�
��6x	p_��x��f�mj�3��b��X�M�H�����WUQ�������m�|�O�rz�0���M��֖8����<�ث�t���3�����\�g���A �^�SlT�Ճ�]���m�-���F�3t>T4�+6�:�/�m���,]GM���˯�����_vC��.�ר'bt�]��Y�	��;��8�Ğ�p��0e�j����;��kA3k�a�@��s|�mrX�a�Þ��2�R%	X�l�aÝ�e���k�o�K�q��V�,�s8G����>Oi��ba4p�I����!��8
(��p��;Jz�����]j-�6��N��gm��9����Ts��>�˨M���������^R�`]]4Z0?y?ş�(��=��HU6���(w�e�������_���<���0���z��ǀ�#�-yɣ`�F����JU\��ه�Mw�c�{���Sa���'� -���@MHiZR��N��A����H"��[k�8$��v�
������<��7�$+3#(�e��H�U�J�}ϥ� ��)7!�0_b&��+5����cy�U��"ZXR��֘-Xqо3���LP'�9�$p +�]� �f��xp�^��%Xh`�)�.,�%�' ����ʑ6��t*
��}Y�\P�w���}��J��`?�a0u;�݈�E��u>��ú_P9wg��z��J�~��4��i[ē��{`����*�_�}�%F�;�{r���F��	�u�������5wlTrG�I;�h.	}Ja�d����Q�#|��s�N�lې���
�v�b��kZQ'x�i������pJ7A�s�~�$�{��Z��Y��|��|WWP߈ A�-k��g;�~�f8m�&�j���Րf��=����p�����bL8ܱ��l�_�pS��X���-�~�8�Yf
P��VS�a�9-�5���J�焗(q�t�J�wq���~�u�g� vw���c�6�J\GE�dӺq8��Ǭ� ��Wb��](�Y�,I����ꦞw�dj9� ~���_^Z}����+��)2�7񕢹���J`8B,�[�ym9��S��#�"��5��Z����V�2o�)[�A��q�k$���?9+�x���-Ԭ]^KE4�P�np��&<�V�`t������v��ʷ���Q���!2�c�2�2,rexBÎ9�����Y�N�Z�Ow)A��T����oit��F����vPQ�R�~��j�CGC�F :�T�x�1IO���1��<��h�aE��9n�7C�P,5�g(}�j_z�f��a񿚼ft�&��������� ��:}�6K"�g�&�K�A(�Z$03�
�'���wV���1 �{�a2�&��T���T �c��՗I�<A� +?��]�f!�\��XCf,�+�!�5���@1�H>����y?��W@�r������!{e`���ՠ��\z�R��}��7�#�hl��zw7�������R��"����JG���%J�0�K ���o�	s���RƮ��?�]4ݤ�n�
����C~�cѮ#��⹻U=�0o�'�3���۫i|8ux  �|3�)k�t�'�5f�n�Wd�ї�$ML�ޚ�(���L:�]�K��@ٍ�B���m+���_-�A1��H�뇚��&��E����2b:~J���f��r��� ��p�u�@��~�e��=����I��;0�e1�� ����#@��ܲ��Fm��y�T�.^���fFNZ��4��P��dmͫr��W%$#����+.֩'x�,���g^�zfp��.h��E�@"����	��i�|�Y�o��ײĊ$��ar��j��#- ��v$���RU.:�1#�Ư/js܎��֠��Gc�ؕ�+` �.�L�ߧ1����T.�P�m��b5��k,�2�cD�T3�����I>Xr(�G�Mi���맫j���Z�H@eA�Ʒ�8g8��e�(fT�t%nk��a�6 �V���I����
\S��Қn�)a�>���F�R���@����Ѳt�t<"4��	D��L���2��,3��C�b/6�k��ŇK"k����T�^Y"�`Tn��xj/TY�4��3�ҿ��������칧���&3"��&X����+<1���&��A�]ã"_Ty\>
%�<g�8�Iq�����C[��	�e�q��L����v�lK!u�&�mq���Z��D��r�krwi�g�4���"��j�ox'��� ]���-�Һ*#
\A��JD��`�Za�	Օ.cjLA7���iL��'���W����TTW��\Qz�����Δ��M�s��S��eV�W�A�_a#� ������;U��Ⱥx���������Ӭ�٠���-Tfo��hr�x ��>�o�`{���ۂ�j<3�e�n�� C~��|�H� .��5�F0f�H���u^#���Nb��Al�2�3�6���?�_�B?"�	ح�pPa!~9f\���[�d�����fnPMp�ʈBFM�)�D���{��tpM���kd��(�b�mY���A��իR�����yG�X��I?���&E���f�>Z��燮gO4�!��ã��cfs��6�t8�Y3�9�L��{!9�HT8�ȩ����@��=�bv�3�<��6�civ��ɷ��d��D�'= ��:��ݖ��I�:Vm}Fi�c����fR���w$z)�凛Nco��4Z��ai�0f�l���܁��✿ă��匕�6�S۬ԛ.��$�6���&v#"�Ƙ�a��R�e��Zh�  ��?'�{��*(����O�6�P�ߠ����~Y&�u g>��˭��:����ঀ�[`EAl�1��w(�^���Q�ˊ��Zt�:]TT�|�s\)��+y��șF���d��:.I��
"W-�� ��s20�͗e�,�ڝ���B��h\���+�B��<[PE����>�r�t��]	��&~/���p�����Ӿ�l m����|��vJڰ�˽�e�ڿ��@��+���!�dg�9O9�s���kNւ�`ϟv7��xC�f�p���z7�sB�k/׿v|!2~A,�r�k �Y������R�)��X�Hl}]���ON�P��2�*�')�$D��X�Ke�V�5p�p�53�*����l߆����/��x�==�ҒZD-~��/��]!�\�����f�s=%	���&�O	�I��\�']���s��,�K#�F`��"��z��4�%�g;�"	��V;O]�3JH[�SIev����:�r<��l�wbWf#���{*�'�
�tp�B��r��1�I%<�e�/c����r
@��^���{nn��7�7D�?�o�����R�?�	 ��â�e�Ft�uA���+^��SO�-?��	�K�a)���
���	��%Eg�ꩉQ�!�w���@� �<#�R�%W_��"���l!^}%K\�y��D���4����-�]?'j6��Р�pR_$�h�_��؍D]�d�H���4�A�ʫ�	�_��)�����v��v�H�\hK�����_]1���л!:$w��D�pkR���3��:�dAۈ�*_7ڪ�>�{���oK:�F�f3_�b{1p��DR�����C�|jFW���=�1��� �k]�6i�~^w4e*��hE1%��t
J�R����ַ5��ts�~��h�nE���w�� �x�c哓;3���?���1Ӵd�1W�̽�{}I�2�m&�6���l��
p~B\)9��`,'ґ�<?'Y<F�?��=&�[��X���#�X0�w֋0�O��f����P��^���fh]q2>%v�G� P)���0͈�UƜT%���JE{�=S}:d�>8]4��*�@P�RI�y�}��@��y�V�5n�2��u���;�$��,!m��5���l��m���JN��}�O������\�0��45=�,XlxV64EB    a53d    1bc0nL��q����ԗ9��r�9m���>�&1jY�f�O��}��@+R��z�Rȿ-��q����/N�;IP�oQ>	�J�D
H�x������e����r��-0�Dt�z]l���O�?Dbhc5�#�lj�-�*���$��b{�$xDW�����K�~���G�V D)қ:xT<�XyW�
�����V\%�ɗ1�4n/8t�;�ϕ��bS{��#����k#����	^�����a���2R�a�_9�@���2[������6*i�}>#�����RHZs��{�<���ݼ$*�L�.g��/��z	����y�����t�i10�_��d���"ђ�׋�S��L.F��(���:�+�W�OjltF��Z�m}p���S ��63]7UC����<F���A[�4y�_^B5n��!�1���$V�8�&E��A$�E��<�X���(��/�U�O�bQ�Zy�����q��Srm��yG��T@�s�0sz��#�$������ �4.�-����k�	�ŷꛒO�ڤ��� �?�.I��W�gs8��4�`��D9��Ln8rD�!v�����ñ�mM�A7�h�~0$�F�tE�����z<p6�[�#�`9m�:G��
0�������h�n��W�A��2h���q~�����9(��\^ �_�;�z��������T���-7B���1Cu�9-�2(�#�X�����CT~�|�R~��_guՆPI�l[,A�ƋEx��w]�W,6kdX>����#+ۚo��O�����mU��һ(:ҧ��1�U�>Z��? �����ҭd�R�rw�����(�Ey[5���3-���L�����������}	�Rg���u�K��]�U֫P���E�ީn/D�j -����w;0����Hշ/h$�DoN��,�"�+Փ^n�^K�zy��T�SЭ۳`P6�7��dOJ���ag|j���fPW�]��p�S׳!����AFݱņ��ʈ����dC�����^���%Ґ7~���(��=22��y��
�Ic��C�Lr��!�5�Ze� <���ͦA����rb��7K�I�K���ȄA-�Y��di!��M�ϙE�S�q�寵̓ՉʒЀ�\Ƌ�M`k
Tzz�7��������V$/O���{V"#,�4��S��o����&`��*��CX7߂T����h�8%M��]����@�
��������/m�fz�X�m�N���n���%?P��!}���o}+�#��q��ع�(+ 8��}5�eutu=>�^�� 5|�9�! )��|ճWR�D,�Nkt�r`�e_C�P�Ug��G��8��bX�U�Jt@&Ly3�ٰ�6���q�La�ZJ�c7�S�[.��i�G]N���[�z��eL�d�[��F|:Ϸ���Sg�~y��ܧ�h��"��<���H�(�^v��C����QzΖ���F����'s�5O�$B����\�:ӂ��{F6m�ߪ�P�4Ko|oǟ�d���޺�	!��6�8j�V�c2��*;�̈�Q�F3�!����}d��Q���0e��c��5�%Z�����A��_ �@�߱T�]�Q�*�^=���!��9�Aj(z�]@۟�1PF������0��'$+^�6S��V����3��xJ6�j՝��4�
�`��㭕�-�i-�Kc�!jp�#���usS�����c԰��~�S����x��ѳh�K�P������6�Σ�w�S'�3�%dP;�^�~޾��^��J�,��!\��/�bO;dB1�">��rc����E/�U��WȬ�n�Iu�L���6�������Q��3[�r:�u����ɇ$LӖSL�����J�� (�=��>���M�$��NJye{�ݫ����2�>gq���dy�&+De�)�,,�:�-騥��#����g�=�o��J;���O�����@*�8�|`[�D�"$#�'�F�X.s��75I�(�E���q'�τ3KI�����E���0C��v�|>hC�{�T�sx���[��a;��n�K�� Hb��*Wo�K�����X��,��	�)�\Fg��:��_V2����Ě�*�(s�6
���ӱ���q7�(ʥ���"����#��,��ƻ��sT X��7Qg�$�?l��߰}����I�nj��c���"��M+����Ej� �>/﫿_��Μ%&��g�����..���0=�7Rxjc�8�S�ӆ���>�	�O!wJme�򡞴<b�j>'z��� h By�nL�d�w�]�`�M�?9b��I1V���`B�2v��`����n���1�}�a,�'p� �7u��R%Ѱ�[��~�dG�ட�,�{� ��+�E�/f�,O}�wi��{��v��)ۃ��-�eŽ��7��$3X�JY�f_��t���޴�#��՟�r'��zp!�nHr�E#˳U1���ݷ�l��d�Nzc �L�Jy�6��=��u�L��z�I��2&��V�
d��v��5hmuK������ڼ�^vkB�щ�������I�)����!M�߬��2/xg:f^6^^�w��F����eikk��_B��f�q��4LĢ^�HO;�1%����@S�4,YJ�\���_��b�gq{޹�?��o�2���~�g�n����p�>tZT����)�v��OF'q[�n{�H�R����݂T&�}烈8M���"���N���8N��>��-x�X�L���'��}�x(\��ݠ�O��(?�8۟mS�g%Zs�ϳ�^�0��|��j�.
�@��%���!!t��![�x��#�{ �?K�%��K9��'���9/>r��շ��S��ǘ�����>��15����'f��/�5 ���rU$y��#�����r�� R.3�b��ҶSb���F�g]��H�?v��^OT�d�I�M��B.ͦe/���WW(�y����s��!���1����wrGs�&�veډaN���AmQ���m��ƪ��Is�U�F�؇>*!\|���5XZ@�E�W��� ���|f���pr4;	�p� ����=�qSqR����M�G�ƣ�O�ǀ����;5�Wb�"���8��d�d(g~_��'�i��p��No�{峝�����Ȅ�X��P�Ep�z%K��q%��~��06��Pmί�������Ǫ��$ =���Z��r �F�ݘ0�-�ہ��ܤ��}����"g�H���+1����R,� �;�J��2\���t�����=����	Bf;�]�,��u�V������`��:'>� N�V��&�H�,�豧�?�����)�`Җ~<��g����b��QQ�G��ōB��t�u_(�A{�*� ٮG���]��o.+q��i�^�DGtL&BJ�货V��\��'�(�8I�LRsN���Qw���_Zpj���=���d]Z}6�3�ln�3%�������'�;^��w[��m˖53�E�Y�ku1"�O	��<Ȋ`7��G� ���f���5F�����t��z�K�[�d�V�sS�(��;�F`_}]�v�,�`�]4�0����t]�ǹ�������=P	��th&�giU �8�l�/"�����T�N�:I�t��f�Ӟ�Ȯ`�����A�m:�/��E(ݢ�]�6��k'������q�`w��i�	 �
�c���~e�;c���=���8�����K������jU��թ��P��NT���&y�d�`��I����x�0��Go�ϒ�9\%��;cd"�ţ���d7����`r�P�l1�����:k�+��\o$��<�|)�=/yf]�hB���ޠf9��0��[H�([�H;ԇ&��b���e�a���ȄTR�z�XH�o��1V�)b�ptM)Eޑ�.�_pk��լ�����g&����s��@7`n.��X�;��R�g��J�mCƯ�N�oA ��8v��{W+��R��ێ(�k����Cυ��Cɻ���x3������l����i"Ftp=߱�5�'d.G�lC�B���f�D��"��W;���n�����p��7��L�aņF�Bc�O)҈59�o� � !���}���K���Fvh�(+Z�]�"ҽ�}�?*B͉RF�vN��{U�HLSO��:а�����(l]��'^�D�p��I?��Ӷ��G>*�ZYL����<��ά;���蒦?��/��RF�PM���~�X�O�j#ӟ�u�J��sr�RE{h"{��K��[,Q����O��v�����V����*�J�V�=�A�y`����2����ƂE���S���/b%���m%u�7�������i#�=���f�>I�WZ�J��&$��a�D���qU0�'��$�h�1מ��!<����o��F@�)B�����U�u����@��4�O�Tbb*��&�yH@�$�3����,���:t>�$d�֣�^D�R��J7�!Y�:�Y7}���P� ]]���D�Z���I��T�_F��1M� ק'��pe�L�e3 ��	�M+�]���2�$�,�ɍ���뇗ݸ&��H���|��X8�
Y����Rh���	<�\��I#�X	-����V�"��fM���[�(�Π����k���W�7`֖��#4X�ӷ,=��Z����,�Y�D��թ{C�֚�_�5K]L eip9�z��A�W"@��~�F/�ƆV��Q�VԂ
 �Yk%|uR#~�u��dp�:d���v��Ŀ�A�\�^Nq��~���gE�F����0����9�,�s_I�v�E��!=��q������b8��yH!�(���/�?�C���ra]��3}�y���G�NX=����Vh|U��/Ȓԅt�F�/����/d��/2�Q���6r��uFs]k�Մ��8�XΛYj�D�Ș�KB^�g��y��O�#�U�ğL���~��K�r� v�0UvJT�	.��D�m��5�� 1�!4��A���K�6�b��r_�{����q���l�~����I�ev�s@/��!�}\�j�);��+RgT�ou+͔��ʠH�b���O1ъO�����=Ը�w�	i����ٓ��k���LK��fG2V.0�����'�"��������c��
��/%-HJ�+���[9~���2,UW5����+::/)�xI��$3���ް�v1I���M��-�x�y^���E=$�ǈ��o�i�%)+� >����D��ޞ�=����$����SM��~�eĩ`���� Ѫ��B�a1�w�>��ȧ�̯�j�/�׼O]Yf�^'0��
6��'<�aC1���O���{#Ib/��u����$ǥ���>+)�:O����O��dY�	�i����l������ڕ��yj&r�&_$+9}��ޮ��hZ$!�FQ��D�n�oLíG{@��e!3��Y�Z�2:�����x�tR�&ߺ�/:gU�XM�6���+�e�{�056O��K齢��w� c��t��pWuU0~wL���T�?�N^�p�3�BvZCpP�K�2�M�����;���yRZa�H~���5k*��:	}�v����*��Z/\*�T�|���=o�09��y�U��ʙř[�&�����I��B��"���?�Q��/2u�n�2!��C9�����\;-YĽi˷��&�SjdS�4�{�L��j7�X�
�"f����/t°G��?������.*��ㆨ�%��NgF��|j�Qk)$	�����dMy�
e������9T�H����4�o
(I������jM�7�ś������I��:;�1�!a� \8G�'Ik��i�b�JPط��W���
�ɯg�c��pb�����R�UN�  ��/�8^>v��p`Yo<t�K�M\�r��{5p�t�p���0��{l����_.���Q `�}�h"�t�)��!�[�OLy�.�kM6��k��5��)��(�L��r�L�l喞1J�7��V�r�!����c��SS���� )ky���R�w�[��-j43�,~��/��2
��WʙM�`�D2�Uo�o�aD��;����c��|�`}�KO�^�V���c�宬��l���d7�f�`�~�ֳ��tw]FP"���	Q��Rk�
âEʱN���g%?%y��q��؁^�lf�t-�������WM=�������� 䝻���0(����#���"!�a�4&�G���0������!�&���@$oo����	�t��iޕ����o~�Ä́���y-FsU�1�f�b��^��Dqġ���Wh���P������Clh1�VMI�B8��Y;�Z^��M&D@�Wژ�ӣ+�3�B&�K��U����<�7�A�b�)D�T^��E�H�,���cڊ<��3Þ/"N��!�]>hT����Q��2 ��h�EiI��I�%4ò��3gn8{��ń�/|^'�/m`�Lܙ�|��"���h��h4��bɛe��j	��1Xx��0�9f�/:&�^�ԑC��객�kn�N�«P��,��*���c@<U�Q�����D��N�*U�O.����!5l%��aݔ�ۢ�t�����G������o�.šʣP&L���=�ff���0IV*;���ZS�v*۪�PsJwl��6��.�Y��2�48��\ �-��X� ۓ=L�8]������@F�ϣ�1q0宭ݍ+��/XF�I�p�/�i�lcR�7��w����c�I����A��lbֺ�"Ly���v�/���J�.�.^�dr�o��E��Ԓ��|�:����:;�Xֽ�����?7���2����Mփ,��,��wMA�3�JB�g)m�{@
!pD�?%,:��A&X:��	��iBixJ&�>��)\8�(PwZ�s��Z৭5s_�k��X�-�l(��D���������}�|��`1wK����%(g��s�^�	�jU�ĥ�g���vkY&���fԛ�[I?�����Ҝ�r