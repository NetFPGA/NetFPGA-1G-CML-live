XlxV64EB    336b     cf0�T(X<ӣ���J@����OӾ���I9���I~��!r�-d�#`6J�?���G����¿M�:M�':f�S����(	^Mtuܔq��E�%�ǒK��B�f��o�x�J�M	�i��-��3iU@`�T��,ʙ���%�h�'Ǟ��)���F��NLUܙ�Is�k�W��Ɯb��{j��P���t+�o�ŋ��MR���[���bk��4T���]$�ۨ|���)oHK�Q8��������^}�@�~�c+�����J����V�5<��)y���mӠ���_҃̃Ұx���lDtVZ'�)A�q';b|v&�]�⢈����	�s���4�}7L֫�*��'����4��y��p���㖂�_y(6�����"�����z��l��F!�w�~1������x����(��mfSC������j��o9��`�QY��s��`ހX�,�k��d"@
�2��,0�S��,(�.��a���z��4�,��E�]���ܔ���ʟ~�auL��+ ;��MČ�?u�Q��-�d�C�d~��z]5yر\	��1�,�yX
X@�R4 ��5Ύ1���s��r��#Pvد�ߪ@�BfT:��2����C�N�oR���|���
EC?m鏲�L��
�r��3%���bHsh�"n�~�I��PC6�п�&���E�c@�~k�@s��]a!G�]90�bmr�����i'4�Ik��$W-h*���E{�g�/9pG3>MtF��/����H���M��	�{5(��)`�i���ydՈ`[���}<N�,�4k�և/o~�i+ƈ�,a�z<�l��b<�#�t�(����� 3�Z�;.�T�-���d	�ۄ��5IS�v��.�`��bh+������%�N��Q@R�=�nM 㶠����G�h�[�0�
��B~z����V�k��Oo� �l�7Z��%2���8t��t���r+�*�0�f5��s��>�L�݁{ֽ���s���o��I����T�U�^듴�����m������� �a�˒�f����&`�*M��T�3��E�h4�SU	C�DrN#D^����qeà"2���x������5nnu0&.��tqT���U�D�Z,�G-�0�ڬ_�X|({�tR�X��PR�G�;"V�@	pҲ�c�̙1�^� o�1�����p�̥VG1��?�v����;��u
���>��C�B��\��e������Sj8�A�h!|0�s^bK�n2f�3D>-�L���k�al�������*���m��d���$�w�E]H��Z����En��ɉF�
�z�f������B�j����̜�
0�tE{�Ey�OS뫡pu:o.1|�����H��8��W�4t*1]�����9%=n:��`se����r�Ge8F#�<�ͷީ���Bë��١�!�ͱ�RC���3��� ��׾��C�������'9eV�Dd��`q��e�Q�I��?�SԀ���ݓ���D��8,��E�ۀ;�~����p^ۄ�����B�τ�--����y��ϣ �����d�!��,o��z�����̚�K���fQp�}��*=�����+���t��8�� ��
�U\�)XP��-ضZ��\�7볬:;p�#O(�r����� �5�,J�s��T���G�� �!�&��dL��	0�y��j�ջn���Jv���B!����@ �vi&ӳ�PH)�!��� ��/�wj�c#43 4��pr��X=1w�T������	��q� �����@"
��/�I"�^͡uw� �)�k+}�-^�9W���������y�>n�����c���o�=���s}�b�N>-o[�&o��\� F�iOB��,���N�d�e�e��U�@�����]ֆ���Zrk�GVcWA=ʬ���2�X
1$��LM�L%�D�1���kQ�8�7d�	�Uվ>�l���u�ס�U:Bu ���jZ�{�y���U�R������9[��Y6���_"S�L�0���͎��+��#�;Prk��8��n�J��[O�^az'�p����`���<��ɏ;�*>�Jl�S���:�� v���tBY�:+���^7��L#��>��]q5�S�jR @K��⹨��,����(/���rfS�$)�5 �����؞k�}����ˆ��10�BJ�Y٣zsh�K�7��c^Y����$��t�������cS��-��?eO�TM�TO���f��	#���Ј��=��,H�1.
Vx�nz�����a�"M��'X� W�a�TA�����mo���cr��+K4���ߴ.��^�SGR�%�\�0j���l���6+������B���"8�#3a�d(�G%)?_pFI�*Z4B���w��;J�Gʥ�ăP� ���?����L�T�"�RF�0p�=l�;*�Mjs��$3R�vۀ�4Oi%���NS�� ֿ�%�z���vV���������lȜ�X���4w���ch�%�������� �y7�u��ð���� �'�b�2�����ܷ����>"�+u�H�Kf��-��W��P/b�p�ˣK��Z5�fJ�N@�r�!;��WoԚ��Q�M�V+��+NeA���*gÐ ���������xk+Z�����r ��1��)��1�̭u�wi�=S�J��q�|Ü��:ٌ�~\���Q*a���Q��4��K�|�9�L�l�7��9��VO�ʓ�_���-�t��C���� �	�"�!ك^Kb(�n�+]�NV�TN��mrDZ�:�͘��LH�>՟{_�Q�Sw*�0���V.Q���${�=��Su�a���/a�1����Ww���D�s���[���h��&W���z��x��Td��K��!ǃa+��0���}�ko�o��6���S��j�&8��M0od*�Do=P���y�7�#�����gp`H"����u�9�QP�]��o�_C��E@n��Q��x�G=3��4<��%�Wk��Z��Ss�v/w�Nh����%��J�@=�f��D�ۣl��T�-�7D% ��e�2���I�J9�Z}Hp�sK�|���A~j�z���= ��T��0���
��!�jS�d�â14ϧJҪH3�;�dW�_h�����VQq��=�t�u��̹��X��dٱ�ve��W���I�6n�M� $���+\Q��6E
`