XlxV64EB    15d6     820��ј!*25ŷ���`�i����SQE<:UfNB�Y�����������t�����ĥ�`W����O�����Z�FV�;��^$x�@���CL�a0�K?uY��]�������Q��L�O����BL���y�Lx�R���tO��.��Ж�uDh�C�A�İk����Zr���ֆ0�e�[��v��+��(Q.�����.��Et_|;FR�X`T=n��h�[@�����d_T־ù�U�0�'gB3�5U�,}�Qc	�o.@��,�i��D��(�4$������*24�f_�	�A���XU��f�`��7C �N�gB��rٰ��cI$�Q�K��U�\�Z4� t��>{�z��J�k5B쿦�T^�{=K�򚎐�ŌZ1�B�xBʋ�˪�ҩM[�9`ϝ���]�i���3`�`l�c3���A&e��a�s��v+�12�wDa�׹ୖ���M�V�;��G\�.jd�빂ߩ�b�fq��|6��Zb�%�餺��ê��E�������9����Q����wM�5�2�θ����E��t��R��K�o�b9�m��������w <��O��Ȝ�m��(�t����´�E�i��k1呶ĵ;[�V=<��������"���U�ˉ�����2]Tw�+6D���{�+���2+�FO��f��D�BPn{C�)�ѐ23��X�	��b{K����(T�|�oc����z#Iq ͮ$j�im>&ՍC5�_��]� 7E�I�ܭ�&�z2���u��)g.[�1h�&R��W��0N�	��QB)&��'Ӡo&�s�q~Y��\�>c��w��حM�-�<������犘�k;���bU�mӁ����G��n�Q�X�6��c�@�����m���9��F֗�'� �Y&�se���, 46�(�*$s?�ۡP����%�"K*͉)Cf���* ������F��X5G�Ƥr�	�}^�9����|=��q_r\S0�>�&�8ݤ� �;����6��M�*Sbm�D~DiMp��j�)ʁ׮TK�K%f7�Ko懊d��)�;J�H��BV+��$�$|�HB�8�ڒ��v��,b�����%��J���F��r8���d���"���O��ߠ9S����3-���¬���$pM�Ä/���q��. 2|~�h+�_uw3QNv���WQL��ڪ�]Z��)b:�c�_
����P)�-_Z�u��e��8�b��L�iV�H�9)�I���zd�t�\�,��]����&�b��}-��I�j:�(�X�C�p���9:��$�9Ԥ�;�,0�4�+y�zjp�I��ުq
�SL�E_� N&�;�w��7�  ����N��L
=M���#�"R�̵��\8d�T�rL\d����:����7��c�g�8m��.k"���:�U�.|h8\c�>]�~�ŉ�VWc���G�qÈi��4U�W�n����.�,��u�0x`e��Zw��G��?�E��?L�~��k��U�����"s���n�8.a߉jK��,�+D��Z18��r�?Y��>ǽ���C3D���4>�L�dd�A���9������ô���"�awDe��<�����Č��V��,RB`�y��zx\�A�J&Q��~%B�o���t�e�� }�|�I��s}zm��<���oG���K�9�r��{�֯&��n�Ã ǜþJ�w�T�2�B���}�R^O��O#%W@@$;Ag��>��Nȅ�b��ϛX�?��g��7t�D6dG?��@�6�ʶ�:%�6)/�-�tnG6NU�Ɉh�)�ڿ)�ZI��s�S�El�H�l��4];2?�ռ�*�U2���}W^�US�+��\�8#���@c�=����]�U�T�$#�`2�79�e@�U~�x73��u!"��A��|}�c@��Uz�.�@1�O��X������]���&�b�Y��%=-^��L�;�q
�jk!��P������]��G5�$��ʁ�b��5\2�:\H��$�u2�@4=��r��O�+%u���`:atS�����%�C�5m��\���F�S8�Ҁ����