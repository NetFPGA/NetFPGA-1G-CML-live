XlxV64EB    566a    1390b��8�-��|IG+��I���t���('���9���`� |la�H�;Ap�G:��ݯ�&r����n?D�`-ųt����`{�j����F��5����m��BK��m?�̳,6�Ǩ�v|���9$z��R�y(��m=�}x�.�	�s�7���'�u�-��)@��ª:躜�r9�ġ��=�5 ��P����Q���V%5V#����{rO&qH�� [%8�{�J���q�(sߔ?��a�΍@n��0���,�>�s_�I0fՖ��:�x3s�_��9�5b~�g`%5�&�WY]���G����!�L�����M�оrw�uvQ dl Uq���Q���V���򀗩3���Jf}7=�9�����S���[��ڎС�Ab�2Svj�N����W�ڂi���6��7���nxD��������\�e�Y�
3�*~���1dan���y�At7���?~D��=�rg��H�(	�}�����4Q���P�Q6�7�M�&�H���A�lBmW��1�<ӓ\��F��ZO��s��vJ�'��,e�VV���X�i�#�^� �?������� �����>В�<�w�pŅ�ʌ.�'D��<W+|�YO9�6O�#f	�* ��jʣt{u �K>Lr_�ϵGC�!�tA�����$.h�_�U	��C8���aqG	����� T���Gx��꫉T���&��6RY6�L�+K��ڤ��$]�ĳ� ԘJj�.����_��U� �m�?���_1s��K���2���pyT��Z��J�F��)cu�`�����Q^��6��N�:�Ա�&�Km9{�a`�,`�Ǿy��j��A���\b>��s߻�E�H��y�|RHg.�Z0�f��?�)��W?%���9��pg�*�s*���6�ސ�i�J4�k��0lq�O�b"��&��/��=sI
�_��ѯ]�$ �+��ٷ��,��c.�#~�V�@OiĨ�sSJ�?��%ɺ��Z<�H�:�@*@y��Wdt�-f��-�,0A℥��0FJ�>vS�(�p!�C��r�u�=x��Z�(��c'�aI(mJ*�U6�B޾��E8��Н;T���y�JY�[��p,�7�>X?��Î#�X����ޞ	94�_��1
�$<�]�^1�q��L�N��Ĳ����ޠ��Q���P�qÿ!��4�5���z���h'���YwW�)9À���SYu�:>O�����^����{i��<����X"�o��l����k�ɽ�W�9A����גev�ӳM�2��f�:������,m0n2���C��RsY���� e�R�W�O�=.O����h4�:Z����J�ޣ4�	ŀ7�T��A�e����.�������F�F��LY/�[���nX����2ij����0<_�S�q�����F��zt�7X]ހ~��&׾H`�Ш�/C,�_�O-�6�gu������L�UF��Pk��g��nL�1�{�O���iI�͎F�yL���R�>��;�u��|ͬr�LDύ�*	�
Qe�^��ܩu��Y
�T��>io��~���<Z���;-QbB�,��}��ڣ���e*55��3����w��S���N��ko��œ���f�T:{�N�O+����$Ǎ�=y-��7%y���K�M��d���"��x�'R/�����r,d,5I{�ZCc �n�7���H����m��z�lҪ� ��!� �Z�����8�=F�y?���((��x�����a��SF�1#'�0o:�|�:ö"(fZh_��8r��j��-�2����JQY>��l��j����FgAR�n`�������$�8��NDrdU{�OC����͛P�AѤ�Ca`ԯ��L�`��J=�O#�o��.A���;$1� ��!�v.%��ux��ӣ��S\�f�8f��,�4����e��Δ��H�W�8I�X5�R��YȤ:�'v�>��9���M; ����q�l.]��x�C�5�������i���)n��Q����5h��:K)�*^����сR��͓��L(ͅ6�Q�I�sQۥ��6hc�C�=J摊���K=(m��7��^�����'����+.��f~&�I���n�`ѡM��sGt��{v�{_�s�Z��q��j�ʓ���/��$�~S��{.D��4�В��@B�Q>(���������&�n��9��hN�6 �baP�Xv�C��%4Ɩ�VG�Ƿ B�PuB�d ��ͷ����)�
����� ]:b��m,[�1Mz���L&A�@̀�|����y���X�o��R�f�ֶ\�;�����1�R���^����
y5��tnw+�=(����P.��-��Z�^U��]�%{�\����n�/0I��=��w�� 05���#�fG���G��}�
�]�.�cck'P.ŹJ�v�";�\���P��X-f� M<����Ř�m��ٶxAؐS��1��\�_	�����\	��U�A�6�rqZȠ�B)��Z������O�]�A��=�A;�HI���w7�WUB=��/$r�~W����8䫁��ڴs3K���Q�:H��̫�\�~�N�++G���mS�7�q��PVD:��AT��{�P~�M��󱽌���vc�bV}�1�{77/C��gV�����s��>�.Bx��f�3P�R��p\�i&�5d�|�`ofZI�K��HF|�(O�8��7�-�s�xBi�M���z�;	l���l�#e-�����[;�z�7Zp�����C�(p��<P�!���ovh�6���3 ��b�@��
2�f�9pT�{��.&�1�q9R�ɓ�$�Jx�;��rN���h-���]�ܙ#h�L`ǕLG��@�5�L�l����2����>A���L\���urѝQ��~��&g���Ίi�Ϳ�%�.u8B�鞯��1��},+�z��zu݈ro�RI�6�OǾ��bO]Gs)7lڈ���[�;�
�fs7hz:{�� �!���^ӯ!(Q�-�b��,0/�1aK�+�=��&��$���4���lV��LQ�)��$�4W��:��-��������C�m����1p�%F�+sN^fK�1S�9��T�"9�+I�}�~σx�}�-1�+��	L�Cā�4�qB�ԥ����>����N�W�h��AUҫ��p<آ��pT��`{v',�

�Ek\(\��4��r�S�t�Ȣ^��Fw�@�o-�y���kZ�V��h,�u�
�����P�Ό��fP��v�S>� \�����5p&�|HF�N/l�^�$-�@�]C!�9����ssȹ��v��θ�*��-)�,�opqN(���#"Y�hwLh���ʳ*c?jt���������ָ��,��|xn�nRyy>�D�# ��7e߀��{Ce3�-���>�	�=�`a�����]jBEԛm�������[%��Q>*��������"�YbM�;h5s��˝yܲ�r��"��z<���k�/�Y�t_�q/%e}���/':�6j����Ы�h��z
���q� %g.�.*��k��[Ӈ[��t�ۆW�Y��A�Se��W�,2t�8��&�Ǫk�1ȴ�9u�"C<Z� �D2���G��N:U�F�ί��_�F��>�j�r<�_� v��9O��e?,�����Qp��������fQ�乚B��{��Xq�?����( �X�I�����!��LdP.�%��> �gN�-݀�0��o&E/arj�L�da��l��ɱ��c��"WZ�%���=it�?�/W��?vη��ttK���4?��if0�5�����$l�+�+eΤt)����*Q=h�(��%Y��<���s,ଗ��oKC��a!��n�Ϋ���[��Vs��V��'3Gv|pWyÌ���ڋ���KK�V�h�4O��%a��]��bT��$�:V��q��|S�� G��`w����h��b�m�2�z���L**G�HG$E��z�M����/Vr���dxw�3.z�$}�J��y&J仺������(�g��MhxI�XG�az��7[5Ҕ��I+.&��mG ��s�v�! �J}Ƞ?#���c�8��h$B� D!���Z��2 ,�0БX���S�?2xM��Ų�ŗ�4��t��SE��n� C�������k�gG(aZ؞�+��:%/��2*�z3fL�CU�쯽����%fR��+�m�(�؃���t�� �9ໂ�����1ޙ]���[c�<%X^F� ��jK�%�5�c@�|J���QU!!�q,V���⮦���Aa=�����x�J�)aφB�U��3���2�CM�T#�Q�K�wh��-��~���������b��,zܫW��//����7'�#� ��i\ր���&�N��E�9�����</�D����- \Z�8�f�,�J�ɷ�M3�ڏT*\:����[�>�	�I�������_�(����4v�Qj�+lStf���LLP��� �.�?��]�=[m5�".����(xq=#�|0&�jۉ������L�[d�(��v��xZ�����#��J�w�@ݰ���Q�1����!�f�'7J*G�OQ8*�$>���c��R��Թ[W���:�a�v�i��\E_�/�����H]�p֍oM����05����J$d�|���k@f��2c���̈́B��Br��TV��R�?R�aG���YW3���PM~"���H5-0ؙ۱�?#Ӈ:����۽�ǜ��<.�M$��!��d�Jv�*�J	P�cJ��0�jB� �T��H�Gj��ŷ�^��_�h����
rQ��Ht���!{[��wYd��b�q��S�]���ƃ�'ߴ�&"���&�'�Y\Ӕ��Po�h3�h�0l�\jf��s"1